/* 
 * EE371 22SP Lab 5 - fancy_animation.sv, May 18, 2022
 * Authors: Haosen Li, Peter Tran
 *
 * Task #3 -- Animation
 *
 * Top level module for line_drawer.sv and clear_screen.sv,
 * creates an animation using the two modules.
 * 
 */
module fancy_animation(input  logic clk, reset,
                 output logic done, color,
                 output logic [10:0] x, y);

    // 26'd50000000 represents 1 second of delay
    logic [25:0] delay_counter;
	logic [7:0] frame_counter;
	logic [7:0] lines_counter;
    logic frame_complete, reset_start;
    // inputs to submodules, manipulate these values
    logic [10:0] x0, y0, x1, y1;
    logic lines_start, clear_start;
    // outputs from submodules, no need to manipulate
    logic [10:0] lines_x, lines_y, clear_x, clear_y;
    logic lines_done, clear_done;

    // instantiate modules
    line_drawer lines(.x(lines_x), .y(lines_y), .reset(lines_start), .done(lines_done), .*);
    clear_screen clear(.x(clear_x), .y(clear_y), .reset(clear_start), .done(clear_done), .*);
    trigger_fsm r_trigger(.in(reset), .out(reset_start), .*);

    // x & y outputs depends on pixel color
    assign x = (color == 1'd1) ? lines_x : clear_x;
    assign y = (color == 1'd1) ? lines_y : clear_y;
    // forever animate? time-based?
    assign done = 1'd0;
    
    always_ff @(posedge clk) begin
        // reset registers
        if (reset) begin
            frame_complete <= 1'd0;
            delay_counter <= 26'd0;
			frame_counter <= 7'd0;
			lines_counter <= 7'd0;
            color <= 1'd0; // black
            x0 <= 11'd0;
            y0 <= 11'd0;
            x1 <= 11'd0;
            y1 <= 11'd0;
        end
        
        if (reset_start) begin
            lines_start <= 1'd1;
            clear_start <= 1'd1;
        end

        // ensures the start signals are only on for one cycle
        if (lines_start == 1'b1)
            lines_start <= 1'b0;
        if (clear_start == 1'b1)
            clear_start <= 1'b0;

        
        /* === FRAMES PER SECOND CONTROL === */

        if (~reset) begin
            // frame delay logic
			if (delay_counter == 26'd5000000) begin
                // increment counters after delay
				if (frame_counter == 7'd111)
					frame_counter <= 7'd0;
				else
					frame_counter <= frame_counter + 1'd1;
                frame_complete <= 1'd0;
                delay_counter <= 26'd0;
                // clear drawing every 1 second
                clear_start <= 1'd1;
                color <= 1'd0; // black
            end else
                // increment delay counter
                delay_counter <= delay_counter + 26'd1;
        end


		/* === ANIMATION FRAMES === */

		// frame 0
		if (frame_counter == 7'd0 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (0, 0) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (0, 0) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (0, 0) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (0, 0) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (0, 0) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (0, 0) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (0, 0) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (0, 0) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (0, 0) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (0, 0) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (0, 0) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (0, 0) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (0, 0) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (0, 0) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (0, 0) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (0, 0) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (0, 0) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (0, 0) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (0, 0) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (0, 0) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (0, 0) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (0, 0) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (0, 0) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (0, 0) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (0, 0) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (0, 0) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (0, 0) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (0, 0) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (0, 0) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (0, 0) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (0, 0) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (0, 0) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (0, 0) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (0, 0) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (0, 0) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (0, 0) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (0, 0) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (0, 0) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (0, 0) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (0, 0) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (0, 0) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (0, 0) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (0, 0) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (0, 0) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (0, 0) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (0, 0) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (0, 0) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (0, 0) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (0, 0) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (0, 0) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (0, 0) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (0, 0) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (0, 0) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (0, 0) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (0, 0) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (0, 0) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (0, 0) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (0, 0) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (0, 0) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (0, 0) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (0, 0) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (0, 0) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (0, 0) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (0, 0) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (0, 0) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (0, 0) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (0, 0) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (0, 0) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (0, 0) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (0, 0) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (0, 0) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (0, 0) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (0, 0) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (0, 0) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (0, 0) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (0, 0) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (0, 0) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (0, 0) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (0, 0) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (0, 0) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (0, 0) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (0, 0) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (0, 0) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (0, 0) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (0, 0) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (0, 0) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (0, 0) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (0, 0) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (0, 0) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (0, 0) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (0, 0) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (0, 0) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (0, 0) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (0, 0) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (0, 0) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (0, 0) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (0, 0) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (0, 0) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (0, 0) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (0, 0) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (0, 0) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (0, 0) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (0, 0) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (0, 0) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (0, 0) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (0, 0) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (0, 0) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (0, 0) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (0, 0) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (0, 0) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (0, 0) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (0, 0) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 1
		if (frame_counter == 7'd1 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (20, 0) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (20, 0) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (20, 0) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (20, 0) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (20, 0) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (20, 0) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (20, 0) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (20, 0) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (20, 0) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (20, 0) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (20, 0) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (20, 0) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (20, 0) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (20, 0) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (20, 0) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (20, 0) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (20, 0) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (20, 0) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (20, 0) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (20, 0) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (20, 0) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (20, 0) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (20, 0) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (20, 0) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (20, 0) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (20, 0) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (20, 0) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (20, 0) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (20, 0) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (20, 0) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (20, 0) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (20, 0) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (20, 0) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (20, 0) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (20, 0) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (20, 0) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (20, 0) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (20, 0) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (20, 0) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (20, 0) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (20, 0) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (20, 0) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (20, 0) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (20, 0) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (20, 0) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (20, 0) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (20, 0) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (20, 0) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (20, 0) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (20, 0) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (20, 0) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (20, 0) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (20, 0) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (20, 0) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (20, 0) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (20, 0) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (20, 0) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (20, 0) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (20, 0) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (20, 0) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (20, 0) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (20, 0) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (20, 0) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (20, 0) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (20, 0) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (20, 0) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (20, 0) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (20, 0) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (20, 0) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (20, 0) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (20, 0) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (20, 0) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (20, 0) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (20, 0) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (20, 0) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (20, 0) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (20, 0) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (20, 0) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (20, 0) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (20, 0) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (20, 0) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (20, 0) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (20, 0) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (20, 0) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (20, 0) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (20, 0) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (20, 0) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (20, 0) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (20, 0) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (20, 0) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (20, 0) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (20, 0) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (20, 0) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (20, 0) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (20, 0) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (20, 0) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (20, 0) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (20, 0) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (20, 0) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (20, 0) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (20, 0) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (20, 0) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (20, 0) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (20, 0) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (20, 0) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (20, 0) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (20, 0) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (20, 0) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (20, 0) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (20, 0) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (20, 0) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (20, 0) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 2
		if (frame_counter == 7'd2 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (40, 0) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (40, 0) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (40, 0) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (40, 0) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (40, 0) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (40, 0) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (40, 0) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (40, 0) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (40, 0) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (40, 0) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (40, 0) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (40, 0) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (40, 0) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (40, 0) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (40, 0) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (40, 0) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (40, 0) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (40, 0) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (40, 0) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (40, 0) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (40, 0) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (40, 0) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (40, 0) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (40, 0) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (40, 0) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (40, 0) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (40, 0) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (40, 0) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (40, 0) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (40, 0) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (40, 0) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (40, 0) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (40, 0) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (40, 0) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (40, 0) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (40, 0) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (40, 0) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (40, 0) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (40, 0) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (40, 0) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (40, 0) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (40, 0) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (40, 0) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (40, 0) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (40, 0) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (40, 0) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (40, 0) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (40, 0) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (40, 0) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (40, 0) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (40, 0) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (40, 0) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (40, 0) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (40, 0) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (40, 0) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (40, 0) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (40, 0) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (40, 0) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (40, 0) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (40, 0) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (40, 0) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (40, 0) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (40, 0) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (40, 0) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (40, 0) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (40, 0) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (40, 0) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (40, 0) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (40, 0) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (40, 0) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (40, 0) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (40, 0) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (40, 0) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (40, 0) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (40, 0) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (40, 0) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (40, 0) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (40, 0) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (40, 0) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (40, 0) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (40, 0) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (40, 0) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (40, 0) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (40, 0) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (40, 0) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (40, 0) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (40, 0) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (40, 0) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (40, 0) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (40, 0) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (40, 0) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (40, 0) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (40, 0) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (40, 0) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (40, 0) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (40, 0) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (40, 0) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (40, 0) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (40, 0) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (40, 0) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (40, 0) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (40, 0) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (40, 0) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (40, 0) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (40, 0) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (40, 0) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (40, 0) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (40, 0) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (40, 0) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (40, 0) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (40, 0) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (40, 0) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 3
		if (frame_counter == 7'd3 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (60, 0) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (60, 0) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (60, 0) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (60, 0) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (60, 0) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (60, 0) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (60, 0) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (60, 0) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (60, 0) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (60, 0) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (60, 0) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (60, 0) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (60, 0) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (60, 0) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (60, 0) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (60, 0) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (60, 0) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (60, 0) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (60, 0) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (60, 0) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (60, 0) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (60, 0) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (60, 0) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (60, 0) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (60, 0) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (60, 0) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (60, 0) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (60, 0) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (60, 0) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (60, 0) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (60, 0) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (60, 0) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (60, 0) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (60, 0) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (60, 0) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (60, 0) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (60, 0) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (60, 0) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (60, 0) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (60, 0) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (60, 0) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (60, 0) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (60, 0) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (60, 0) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (60, 0) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (60, 0) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (60, 0) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (60, 0) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (60, 0) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (60, 0) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (60, 0) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (60, 0) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (60, 0) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (60, 0) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (60, 0) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (60, 0) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (60, 0) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (60, 0) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (60, 0) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (60, 0) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (60, 0) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (60, 0) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (60, 0) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (60, 0) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (60, 0) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (60, 0) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (60, 0) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (60, 0) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (60, 0) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (60, 0) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (60, 0) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (60, 0) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (60, 0) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (60, 0) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (60, 0) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (60, 0) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (60, 0) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (60, 0) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (60, 0) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (60, 0) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (60, 0) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (60, 0) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (60, 0) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (60, 0) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (60, 0) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (60, 0) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (60, 0) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (60, 0) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (60, 0) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (60, 0) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (60, 0) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (60, 0) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (60, 0) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (60, 0) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (60, 0) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (60, 0) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (60, 0) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (60, 0) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (60, 0) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (60, 0) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (60, 0) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (60, 0) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (60, 0) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (60, 0) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (60, 0) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (60, 0) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (60, 0) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (60, 0) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (60, 0) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (60, 0) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (60, 0) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (60, 0) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 4
		if (frame_counter == 7'd4 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (80, 0) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (80, 0) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (80, 0) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (80, 0) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (80, 0) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (80, 0) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (80, 0) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (80, 0) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (80, 0) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (80, 0) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (80, 0) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (80, 0) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (80, 0) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (80, 0) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (80, 0) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (80, 0) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (80, 0) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (80, 0) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (80, 0) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (80, 0) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (80, 0) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (80, 0) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (80, 0) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (80, 0) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (80, 0) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (80, 0) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (80, 0) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (80, 0) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (80, 0) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (80, 0) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (80, 0) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (80, 0) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (80, 0) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (80, 0) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (80, 0) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (80, 0) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (80, 0) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (80, 0) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (80, 0) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (80, 0) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (80, 0) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (80, 0) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (80, 0) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (80, 0) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (80, 0) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (80, 0) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (80, 0) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (80, 0) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (80, 0) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (80, 0) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (80, 0) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (80, 0) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (80, 0) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (80, 0) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (80, 0) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (80, 0) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (80, 0) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (80, 0) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (80, 0) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (80, 0) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (80, 0) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (80, 0) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (80, 0) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (80, 0) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (80, 0) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (80, 0) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (80, 0) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (80, 0) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (80, 0) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (80, 0) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (80, 0) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (80, 0) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (80, 0) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (80, 0) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (80, 0) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (80, 0) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (80, 0) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (80, 0) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (80, 0) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (80, 0) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (80, 0) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (80, 0) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (80, 0) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (80, 0) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (80, 0) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (80, 0) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (80, 0) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (80, 0) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (80, 0) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (80, 0) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (80, 0) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (80, 0) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (80, 0) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (80, 0) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (80, 0) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (80, 0) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (80, 0) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (80, 0) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (80, 0) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (80, 0) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (80, 0) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (80, 0) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (80, 0) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (80, 0) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (80, 0) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (80, 0) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (80, 0) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (80, 0) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (80, 0) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (80, 0) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (80, 0) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (80, 0) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 5
		if (frame_counter == 7'd5 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (100, 0) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (100, 0) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (100, 0) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (100, 0) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (100, 0) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (100, 0) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (100, 0) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (100, 0) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (100, 0) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (100, 0) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (100, 0) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (100, 0) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (100, 0) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (100, 0) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (100, 0) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (100, 0) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (100, 0) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (100, 0) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (100, 0) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (100, 0) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (100, 0) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (100, 0) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (100, 0) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (100, 0) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (100, 0) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (100, 0) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (100, 0) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (100, 0) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (100, 0) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (100, 0) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (100, 0) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (100, 0) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (100, 0) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (100, 0) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (100, 0) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (100, 0) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (100, 0) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (100, 0) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (100, 0) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (100, 0) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (100, 0) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (100, 0) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (100, 0) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (100, 0) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (100, 0) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (100, 0) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (100, 0) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (100, 0) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (100, 0) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (100, 0) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (100, 0) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (100, 0) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (100, 0) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (100, 0) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (100, 0) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (100, 0) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (100, 0) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (100, 0) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (100, 0) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (100, 0) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (100, 0) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (100, 0) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (100, 0) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (100, 0) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (100, 0) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (100, 0) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (100, 0) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (100, 0) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (100, 0) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (100, 0) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (100, 0) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (100, 0) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (100, 0) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (100, 0) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (100, 0) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (100, 0) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (100, 0) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (100, 0) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (100, 0) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (100, 0) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (100, 0) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (100, 0) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (100, 0) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (100, 0) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (100, 0) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (100, 0) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (100, 0) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (100, 0) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (100, 0) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (100, 0) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (100, 0) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (100, 0) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (100, 0) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (100, 0) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (100, 0) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (100, 0) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (100, 0) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (100, 0) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (100, 0) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (100, 0) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (100, 0) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (100, 0) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (100, 0) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (100, 0) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (100, 0) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (100, 0) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (100, 0) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (100, 0) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (100, 0) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (100, 0) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (100, 0) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (100, 0) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 6
		if (frame_counter == 7'd6 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (120, 0) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (120, 0) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (120, 0) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (120, 0) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (120, 0) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (120, 0) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (120, 0) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (120, 0) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (120, 0) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (120, 0) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (120, 0) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (120, 0) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (120, 0) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (120, 0) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (120, 0) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (120, 0) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (120, 0) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (120, 0) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (120, 0) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (120, 0) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (120, 0) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (120, 0) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (120, 0) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (120, 0) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (120, 0) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (120, 0) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (120, 0) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (120, 0) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (120, 0) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (120, 0) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (120, 0) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (120, 0) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (120, 0) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (120, 0) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (120, 0) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (120, 0) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (120, 0) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (120, 0) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (120, 0) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (120, 0) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (120, 0) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (120, 0) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (120, 0) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (120, 0) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (120, 0) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (120, 0) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (120, 0) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (120, 0) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (120, 0) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (120, 0) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (120, 0) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (120, 0) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (120, 0) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (120, 0) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (120, 0) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (120, 0) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (120, 0) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (120, 0) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (120, 0) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (120, 0) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (120, 0) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (120, 0) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (120, 0) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (120, 0) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (120, 0) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (120, 0) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (120, 0) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (120, 0) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (120, 0) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (120, 0) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (120, 0) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (120, 0) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (120, 0) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (120, 0) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (120, 0) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (120, 0) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (120, 0) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (120, 0) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (120, 0) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (120, 0) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (120, 0) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (120, 0) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (120, 0) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (120, 0) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (120, 0) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (120, 0) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (120, 0) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (120, 0) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (120, 0) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (120, 0) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (120, 0) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (120, 0) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (120, 0) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (120, 0) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (120, 0) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (120, 0) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (120, 0) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (120, 0) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (120, 0) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (120, 0) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (120, 0) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (120, 0) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (120, 0) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (120, 0) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (120, 0) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (120, 0) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (120, 0) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (120, 0) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (120, 0) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (120, 0) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (120, 0) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (120, 0) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 7
		if (frame_counter == 7'd7 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (140, 0) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (140, 0) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (140, 0) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (140, 0) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (140, 0) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (140, 0) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (140, 0) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (140, 0) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (140, 0) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (140, 0) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (140, 0) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (140, 0) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (140, 0) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (140, 0) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (140, 0) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (140, 0) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (140, 0) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (140, 0) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (140, 0) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (140, 0) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (140, 0) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (140, 0) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (140, 0) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (140, 0) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (140, 0) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (140, 0) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (140, 0) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (140, 0) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (140, 0) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (140, 0) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (140, 0) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (140, 0) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (140, 0) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (140, 0) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (140, 0) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (140, 0) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (140, 0) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (140, 0) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (140, 0) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (140, 0) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (140, 0) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (140, 0) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (140, 0) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (140, 0) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (140, 0) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (140, 0) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (140, 0) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (140, 0) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (140, 0) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (140, 0) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (140, 0) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (140, 0) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (140, 0) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (140, 0) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (140, 0) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (140, 0) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (140, 0) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (140, 0) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (140, 0) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (140, 0) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (140, 0) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (140, 0) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (140, 0) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (140, 0) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (140, 0) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (140, 0) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (140, 0) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (140, 0) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (140, 0) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (140, 0) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (140, 0) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (140, 0) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (140, 0) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (140, 0) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (140, 0) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (140, 0) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (140, 0) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (140, 0) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (140, 0) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (140, 0) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (140, 0) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (140, 0) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (140, 0) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (140, 0) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (140, 0) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (140, 0) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (140, 0) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (140, 0) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (140, 0) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (140, 0) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (140, 0) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (140, 0) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (140, 0) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (140, 0) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (140, 0) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (140, 0) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (140, 0) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (140, 0) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (140, 0) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (140, 0) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (140, 0) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (140, 0) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (140, 0) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (140, 0) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (140, 0) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (140, 0) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (140, 0) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (140, 0) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (140, 0) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (140, 0) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (140, 0) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (140, 0) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 8
		if (frame_counter == 7'd8 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (160, 0) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (160, 0) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (160, 0) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (160, 0) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (160, 0) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (160, 0) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (160, 0) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (160, 0) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (160, 0) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (160, 0) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (160, 0) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (160, 0) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (160, 0) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (160, 0) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (160, 0) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (160, 0) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (160, 0) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (160, 0) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (160, 0) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (160, 0) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (160, 0) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (160, 0) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (160, 0) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (160, 0) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (160, 0) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (160, 0) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (160, 0) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (160, 0) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (160, 0) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (160, 0) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (160, 0) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (160, 0) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (160, 0) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (160, 0) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (160, 0) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (160, 0) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (160, 0) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (160, 0) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (160, 0) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (160, 0) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (160, 0) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (160, 0) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (160, 0) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (160, 0) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (160, 0) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (160, 0) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (160, 0) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (160, 0) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (160, 0) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (160, 0) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (160, 0) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (160, 0) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (160, 0) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (160, 0) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (160, 0) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (160, 0) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (160, 0) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (160, 0) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (160, 0) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (160, 0) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (160, 0) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (160, 0) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (160, 0) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (160, 0) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (160, 0) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (160, 0) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (160, 0) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (160, 0) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (160, 0) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (160, 0) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (160, 0) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (160, 0) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (160, 0) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (160, 0) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (160, 0) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (160, 0) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (160, 0) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (160, 0) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (160, 0) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (160, 0) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (160, 0) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (160, 0) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (160, 0) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (160, 0) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (160, 0) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (160, 0) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (160, 0) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (160, 0) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (160, 0) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (160, 0) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (160, 0) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (160, 0) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (160, 0) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (160, 0) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (160, 0) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (160, 0) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (160, 0) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (160, 0) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (160, 0) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (160, 0) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (160, 0) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (160, 0) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (160, 0) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (160, 0) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (160, 0) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (160, 0) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (160, 0) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (160, 0) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (160, 0) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (160, 0) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (160, 0) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (160, 0) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 9
		if (frame_counter == 7'd9 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (180, 0) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (180, 0) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (180, 0) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (180, 0) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (180, 0) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (180, 0) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (180, 0) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (180, 0) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (180, 0) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (180, 0) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (180, 0) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (180, 0) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (180, 0) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (180, 0) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (180, 0) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (180, 0) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (180, 0) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (180, 0) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (180, 0) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (180, 0) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (180, 0) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (180, 0) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (180, 0) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (180, 0) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (180, 0) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (180, 0) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (180, 0) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (180, 0) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (180, 0) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (180, 0) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (180, 0) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (180, 0) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (180, 0) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (180, 0) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (180, 0) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (180, 0) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (180, 0) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (180, 0) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (180, 0) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (180, 0) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (180, 0) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (180, 0) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (180, 0) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (180, 0) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (180, 0) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (180, 0) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (180, 0) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (180, 0) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (180, 0) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (180, 0) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (180, 0) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (180, 0) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (180, 0) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (180, 0) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (180, 0) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (180, 0) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (180, 0) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (180, 0) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (180, 0) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (180, 0) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (180, 0) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (180, 0) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (180, 0) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (180, 0) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (180, 0) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (180, 0) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (180, 0) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (180, 0) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (180, 0) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (180, 0) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (180, 0) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (180, 0) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (180, 0) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (180, 0) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (180, 0) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (180, 0) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (180, 0) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (180, 0) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (180, 0) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (180, 0) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (180, 0) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (180, 0) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (180, 0) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (180, 0) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (180, 0) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (180, 0) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (180, 0) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (180, 0) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (180, 0) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (180, 0) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (180, 0) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (180, 0) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (180, 0) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (180, 0) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (180, 0) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (180, 0) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (180, 0) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (180, 0) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (180, 0) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (180, 0) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (180, 0) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (180, 0) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (180, 0) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (180, 0) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (180, 0) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (180, 0) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (180, 0) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (180, 0) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (180, 0) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (180, 0) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (180, 0) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (180, 0) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 10
		if (frame_counter == 7'd10 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (200, 0) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (200, 0) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (200, 0) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (200, 0) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (200, 0) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (200, 0) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (200, 0) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (200, 0) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (200, 0) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (200, 0) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (200, 0) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (200, 0) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (200, 0) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (200, 0) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (200, 0) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (200, 0) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (200, 0) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (200, 0) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (200, 0) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (200, 0) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (200, 0) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (200, 0) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (200, 0) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (200, 0) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (200, 0) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (200, 0) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (200, 0) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (200, 0) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (200, 0) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (200, 0) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (200, 0) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (200, 0) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (200, 0) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (200, 0) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (200, 0) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (200, 0) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (200, 0) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (200, 0) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (200, 0) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (200, 0) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (200, 0) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (200, 0) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (200, 0) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (200, 0) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (200, 0) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (200, 0) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (200, 0) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (200, 0) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (200, 0) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (200, 0) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (200, 0) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (200, 0) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (200, 0) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (200, 0) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (200, 0) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (200, 0) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (200, 0) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (200, 0) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (200, 0) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (200, 0) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (200, 0) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (200, 0) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (200, 0) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (200, 0) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (200, 0) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (200, 0) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (200, 0) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (200, 0) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (200, 0) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (200, 0) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (200, 0) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (200, 0) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (200, 0) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (200, 0) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (200, 0) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (200, 0) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (200, 0) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (200, 0) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (200, 0) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (200, 0) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (200, 0) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (200, 0) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (200, 0) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (200, 0) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (200, 0) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (200, 0) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (200, 0) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (200, 0) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (200, 0) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (200, 0) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (200, 0) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (200, 0) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (200, 0) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (200, 0) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (200, 0) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (200, 0) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (200, 0) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (200, 0) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (200, 0) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (200, 0) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (200, 0) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (200, 0) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (200, 0) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (200, 0) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (200, 0) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (200, 0) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (200, 0) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (200, 0) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (200, 0) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (200, 0) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (200, 0) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (200, 0) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 11
		if (frame_counter == 7'd11 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (220, 0) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (220, 0) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (220, 0) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (220, 0) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (220, 0) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (220, 0) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (220, 0) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (220, 0) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (220, 0) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (220, 0) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (220, 0) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (220, 0) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (220, 0) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (220, 0) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (220, 0) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (220, 0) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (220, 0) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (220, 0) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (220, 0) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (220, 0) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (220, 0) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (220, 0) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (220, 0) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (220, 0) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (220, 0) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (220, 0) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (220, 0) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (220, 0) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (220, 0) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (220, 0) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (220, 0) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (220, 0) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (220, 0) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (220, 0) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (220, 0) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (220, 0) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (220, 0) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (220, 0) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (220, 0) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (220, 0) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (220, 0) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (220, 0) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (220, 0) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (220, 0) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (220, 0) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (220, 0) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (220, 0) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (220, 0) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (220, 0) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (220, 0) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (220, 0) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (220, 0) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (220, 0) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (220, 0) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (220, 0) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (220, 0) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (220, 0) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (220, 0) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (220, 0) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (220, 0) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (220, 0) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (220, 0) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (220, 0) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (220, 0) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (220, 0) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (220, 0) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (220, 0) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (220, 0) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (220, 0) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (220, 0) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (220, 0) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (220, 0) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (220, 0) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (220, 0) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (220, 0) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (220, 0) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (220, 0) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (220, 0) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (220, 0) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (220, 0) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (220, 0) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (220, 0) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (220, 0) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (220, 0) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (220, 0) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (220, 0) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (220, 0) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (220, 0) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (220, 0) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (220, 0) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (220, 0) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (220, 0) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (220, 0) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (220, 0) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (220, 0) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (220, 0) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (220, 0) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (220, 0) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (220, 0) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (220, 0) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (220, 0) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (220, 0) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (220, 0) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (220, 0) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (220, 0) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (220, 0) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (220, 0) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (220, 0) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (220, 0) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (220, 0) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (220, 0) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (220, 0) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 12
		if (frame_counter == 7'd12 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (240, 0) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (240, 0) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (240, 0) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (240, 0) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (240, 0) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (240, 0) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (240, 0) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (240, 0) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (240, 0) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (240, 0) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (240, 0) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (240, 0) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (240, 0) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (240, 0) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (240, 0) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (240, 0) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (240, 0) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (240, 0) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (240, 0) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (240, 0) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (240, 0) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (240, 0) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (240, 0) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (240, 0) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (240, 0) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (240, 0) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (240, 0) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (240, 0) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (240, 0) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (240, 0) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (240, 0) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (240, 0) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (240, 0) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (240, 0) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (240, 0) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (240, 0) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (240, 0) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (240, 0) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (240, 0) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (240, 0) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (240, 0) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (240, 0) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (240, 0) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (240, 0) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (240, 0) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (240, 0) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (240, 0) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (240, 0) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (240, 0) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (240, 0) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (240, 0) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (240, 0) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (240, 0) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (240, 0) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (240, 0) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (240, 0) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (240, 0) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (240, 0) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (240, 0) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (240, 0) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (240, 0) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (240, 0) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (240, 0) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (240, 0) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (240, 0) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (240, 0) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (240, 0) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (240, 0) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (240, 0) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (240, 0) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (240, 0) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (240, 0) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (240, 0) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (240, 0) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (240, 0) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (240, 0) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (240, 0) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (240, 0) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (240, 0) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (240, 0) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (240, 0) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (240, 0) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (240, 0) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (240, 0) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (240, 0) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (240, 0) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (240, 0) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (240, 0) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (240, 0) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (240, 0) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (240, 0) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (240, 0) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (240, 0) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (240, 0) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (240, 0) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (240, 0) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (240, 0) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (240, 0) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (240, 0) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (240, 0) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (240, 0) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (240, 0) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (240, 0) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (240, 0) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (240, 0) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (240, 0) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (240, 0) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (240, 0) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (240, 0) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (240, 0) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (240, 0) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (240, 0) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 13
		if (frame_counter == 7'd13 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (260, 0) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (260, 0) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (260, 0) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (260, 0) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (260, 0) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (260, 0) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (260, 0) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (260, 0) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (260, 0) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (260, 0) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (260, 0) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (260, 0) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (260, 0) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (260, 0) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (260, 0) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (260, 0) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (260, 0) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (260, 0) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (260, 0) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (260, 0) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (260, 0) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (260, 0) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (260, 0) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (260, 0) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (260, 0) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (260, 0) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (260, 0) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (260, 0) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (260, 0) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (260, 0) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (260, 0) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (260, 0) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (260, 0) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (260, 0) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (260, 0) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (260, 0) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (260, 0) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (260, 0) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (260, 0) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (260, 0) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (260, 0) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (260, 0) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (260, 0) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (260, 0) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (260, 0) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (260, 0) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (260, 0) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (260, 0) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (260, 0) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (260, 0) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (260, 0) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (260, 0) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (260, 0) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (260, 0) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (260, 0) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (260, 0) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (260, 0) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (260, 0) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (260, 0) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (260, 0) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (260, 0) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (260, 0) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (260, 0) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (260, 0) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (260, 0) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (260, 0) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (260, 0) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (260, 0) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (260, 0) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (260, 0) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (260, 0) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (260, 0) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (260, 0) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (260, 0) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (260, 0) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (260, 0) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (260, 0) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (260, 0) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (260, 0) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (260, 0) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (260, 0) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (260, 0) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (260, 0) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (260, 0) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (260, 0) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (260, 0) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (260, 0) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (260, 0) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (260, 0) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (260, 0) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (260, 0) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (260, 0) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (260, 0) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (260, 0) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (260, 0) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (260, 0) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (260, 0) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (260, 0) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (260, 0) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (260, 0) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (260, 0) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (260, 0) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (260, 0) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (260, 0) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (260, 0) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (260, 0) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (260, 0) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (260, 0) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (260, 0) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (260, 0) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (260, 0) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (260, 0) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 14
		if (frame_counter == 7'd14 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (280, 0) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (280, 0) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (280, 0) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (280, 0) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (280, 0) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (280, 0) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (280, 0) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (280, 0) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (280, 0) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (280, 0) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (280, 0) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (280, 0) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (280, 0) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (280, 0) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (280, 0) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (280, 0) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (280, 0) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (280, 0) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (280, 0) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (280, 0) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (280, 0) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (280, 0) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (280, 0) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (280, 0) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (280, 0) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (280, 0) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (280, 0) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (280, 0) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (280, 0) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (280, 0) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (280, 0) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (280, 0) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (280, 0) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (280, 0) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (280, 0) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (280, 0) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (280, 0) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (280, 0) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (280, 0) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (280, 0) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (280, 0) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (280, 0) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (280, 0) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (280, 0) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (280, 0) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (280, 0) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (280, 0) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (280, 0) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (280, 0) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (280, 0) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (280, 0) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (280, 0) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (280, 0) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (280, 0) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (280, 0) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (280, 0) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (280, 0) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (280, 0) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (280, 0) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (280, 0) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (280, 0) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (280, 0) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (280, 0) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (280, 0) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (280, 0) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (280, 0) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (280, 0) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (280, 0) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (280, 0) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (280, 0) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (280, 0) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (280, 0) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (280, 0) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (280, 0) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (280, 0) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (280, 0) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (280, 0) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (280, 0) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (280, 0) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (280, 0) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (280, 0) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (280, 0) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (280, 0) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (280, 0) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (280, 0) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (280, 0) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (280, 0) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (280, 0) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (280, 0) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (280, 0) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (280, 0) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (280, 0) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (280, 0) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (280, 0) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (280, 0) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (280, 0) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (280, 0) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (280, 0) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (280, 0) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (280, 0) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (280, 0) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (280, 0) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (280, 0) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (280, 0) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (280, 0) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (280, 0) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (280, 0) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (280, 0) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (280, 0) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (280, 0) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (280, 0) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (280, 0) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 15
		if (frame_counter == 7'd15 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (300, 0) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (300, 0) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (300, 0) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (300, 0) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (300, 0) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (300, 0) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (300, 0) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (300, 0) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (300, 0) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (300, 0) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (300, 0) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (300, 0) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (300, 0) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (300, 0) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (300, 0) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (300, 0) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (300, 0) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (300, 0) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (300, 0) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (300, 0) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (300, 0) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (300, 0) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (300, 0) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (300, 0) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (300, 0) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (300, 0) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (300, 0) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (300, 0) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (300, 0) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (300, 0) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (300, 0) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (300, 0) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (300, 0) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (300, 0) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (300, 0) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (300, 0) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (300, 0) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (300, 0) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (300, 0) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (300, 0) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (300, 0) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (300, 0) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (300, 0) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (300, 0) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (300, 0) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (300, 0) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (300, 0) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (300, 0) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (300, 0) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (300, 0) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (300, 0) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (300, 0) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (300, 0) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (300, 0) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (300, 0) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (300, 0) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (300, 0) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (300, 0) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (300, 0) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (300, 0) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (300, 0) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (300, 0) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (300, 0) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (300, 0) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (300, 0) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (300, 0) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (300, 0) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (300, 0) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (300, 0) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (300, 0) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (300, 0) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (300, 0) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (300, 0) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (300, 0) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (300, 0) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (300, 0) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (300, 0) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (300, 0) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (300, 0) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (300, 0) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (300, 0) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (300, 0) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (300, 0) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (300, 0) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (300, 0) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (300, 0) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (300, 0) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (300, 0) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (300, 0) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (300, 0) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (300, 0) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (300, 0) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (300, 0) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (300, 0) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (300, 0) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (300, 0) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (300, 0) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (300, 0) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (300, 0) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (300, 0) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (300, 0) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (300, 0) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (300, 0) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (300, 0) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (300, 0) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (300, 0) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (300, 0) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (300, 0) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (300, 0) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (300, 0) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (300, 0) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (300, 0) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 16
		if (frame_counter == 7'd16 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (320, 0) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (320, 0) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (320, 0) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (320, 0) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (320, 0) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (320, 0) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (320, 0) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (320, 0) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (320, 0) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (320, 0) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (320, 0) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (320, 0) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (320, 0) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (320, 0) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (320, 0) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (320, 0) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (320, 0) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (320, 0) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (320, 0) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (320, 0) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (320, 0) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (320, 0) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (320, 0) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (320, 0) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (320, 0) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (320, 0) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (320, 0) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (320, 0) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (320, 0) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (320, 0) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (320, 0) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (320, 0) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (320, 0) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (320, 0) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (320, 0) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (320, 0) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (320, 0) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (320, 0) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (320, 0) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (320, 0) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (320, 0) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (320, 0) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (320, 0) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (320, 0) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (320, 0) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (320, 0) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (320, 0) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (320, 0) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (320, 0) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (320, 0) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (320, 0) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (320, 0) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (320, 0) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (320, 0) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (320, 0) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (320, 0) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (320, 0) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (320, 0) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (320, 0) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (320, 0) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (320, 0) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (320, 0) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (320, 0) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (320, 0) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (320, 0) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (320, 0) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (320, 0) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (320, 0) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (320, 0) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (320, 0) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (320, 0) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (320, 0) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (320, 0) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (320, 0) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (320, 0) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (320, 0) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (320, 0) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (320, 0) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (320, 0) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (320, 0) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (320, 0) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (320, 0) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (320, 0) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (320, 0) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (320, 0) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (320, 0) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (320, 0) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (320, 0) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (320, 0) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (320, 0) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (320, 0) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (320, 0) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (320, 0) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (320, 0) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (320, 0) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (320, 0) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (320, 0) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (320, 0) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (320, 0) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (320, 0) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (320, 0) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (320, 0) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (320, 0) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (320, 0) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (320, 0) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (320, 0) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (320, 0) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (320, 0) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (320, 0) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (320, 0) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (320, 0) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (320, 0) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 17
		if (frame_counter == 7'd17 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (340, 0) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (340, 0) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (340, 0) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (340, 0) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (340, 0) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (340, 0) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (340, 0) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (340, 0) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (340, 0) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (340, 0) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (340, 0) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (340, 0) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (340, 0) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (340, 0) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (340, 0) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (340, 0) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (340, 0) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (340, 0) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (340, 0) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (340, 0) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (340, 0) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (340, 0) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (340, 0) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (340, 0) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (340, 0) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (340, 0) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (340, 0) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (340, 0) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (340, 0) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (340, 0) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (340, 0) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (340, 0) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (340, 0) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (340, 0) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (340, 0) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (340, 0) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (340, 0) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (340, 0) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (340, 0) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (340, 0) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (340, 0) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (340, 0) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (340, 0) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (340, 0) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (340, 0) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (340, 0) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (340, 0) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (340, 0) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (340, 0) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (340, 0) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (340, 0) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (340, 0) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (340, 0) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (340, 0) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (340, 0) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (340, 0) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (340, 0) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (340, 0) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (340, 0) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (340, 0) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (340, 0) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (340, 0) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (340, 0) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (340, 0) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (340, 0) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (340, 0) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (340, 0) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (340, 0) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (340, 0) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (340, 0) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (340, 0) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (340, 0) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (340, 0) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (340, 0) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (340, 0) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (340, 0) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (340, 0) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (340, 0) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (340, 0) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (340, 0) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (340, 0) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (340, 0) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (340, 0) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (340, 0) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (340, 0) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (340, 0) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (340, 0) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (340, 0) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (340, 0) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (340, 0) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (340, 0) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (340, 0) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (340, 0) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (340, 0) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (340, 0) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (340, 0) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (340, 0) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (340, 0) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (340, 0) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (340, 0) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (340, 0) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (340, 0) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (340, 0) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (340, 0) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (340, 0) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (340, 0) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (340, 0) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (340, 0) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (340, 0) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (340, 0) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (340, 0) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (340, 0) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 18
		if (frame_counter == 7'd18 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (360, 0) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (360, 0) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (360, 0) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (360, 0) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (360, 0) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (360, 0) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (360, 0) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (360, 0) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (360, 0) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (360, 0) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (360, 0) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (360, 0) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (360, 0) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (360, 0) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (360, 0) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (360, 0) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (360, 0) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (360, 0) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (360, 0) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (360, 0) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (360, 0) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (360, 0) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (360, 0) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (360, 0) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (360, 0) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (360, 0) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (360, 0) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (360, 0) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (360, 0) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (360, 0) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (360, 0) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (360, 0) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (360, 0) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (360, 0) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (360, 0) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (360, 0) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (360, 0) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (360, 0) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (360, 0) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (360, 0) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (360, 0) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (360, 0) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (360, 0) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (360, 0) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (360, 0) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (360, 0) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (360, 0) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (360, 0) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (360, 0) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (360, 0) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (360, 0) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (360, 0) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (360, 0) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (360, 0) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (360, 0) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (360, 0) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (360, 0) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (360, 0) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (360, 0) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (360, 0) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (360, 0) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (360, 0) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (360, 0) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (360, 0) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (360, 0) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (360, 0) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (360, 0) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (360, 0) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (360, 0) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (360, 0) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (360, 0) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (360, 0) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (360, 0) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (360, 0) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (360, 0) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (360, 0) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (360, 0) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (360, 0) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (360, 0) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (360, 0) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (360, 0) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (360, 0) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (360, 0) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (360, 0) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (360, 0) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (360, 0) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (360, 0) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (360, 0) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (360, 0) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (360, 0) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (360, 0) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (360, 0) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (360, 0) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (360, 0) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (360, 0) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (360, 0) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (360, 0) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (360, 0) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (360, 0) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (360, 0) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (360, 0) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (360, 0) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (360, 0) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (360, 0) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (360, 0) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (360, 0) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (360, 0) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (360, 0) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (360, 0) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (360, 0) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (360, 0) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (360, 0) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 19
		if (frame_counter == 7'd19 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (380, 0) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (380, 0) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (380, 0) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (380, 0) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (380, 0) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (380, 0) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (380, 0) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (380, 0) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (380, 0) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (380, 0) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (380, 0) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (380, 0) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (380, 0) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (380, 0) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (380, 0) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (380, 0) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (380, 0) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (380, 0) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (380, 0) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (380, 0) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (380, 0) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (380, 0) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (380, 0) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (380, 0) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (380, 0) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (380, 0) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (380, 0) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (380, 0) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (380, 0) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (380, 0) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (380, 0) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (380, 0) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (380, 0) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (380, 0) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (380, 0) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (380, 0) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (380, 0) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (380, 0) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (380, 0) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (380, 0) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (380, 0) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (380, 0) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (380, 0) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (380, 0) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (380, 0) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (380, 0) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (380, 0) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (380, 0) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (380, 0) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (380, 0) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (380, 0) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (380, 0) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (380, 0) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (380, 0) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (380, 0) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (380, 0) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (380, 0) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (380, 0) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (380, 0) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (380, 0) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (380, 0) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (380, 0) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (380, 0) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (380, 0) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (380, 0) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (380, 0) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (380, 0) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (380, 0) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (380, 0) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (380, 0) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (380, 0) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (380, 0) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (380, 0) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (380, 0) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (380, 0) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (380, 0) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (380, 0) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (380, 0) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (380, 0) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (380, 0) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (380, 0) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (380, 0) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (380, 0) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (380, 0) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (380, 0) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (380, 0) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (380, 0) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (380, 0) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (380, 0) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (380, 0) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (380, 0) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (380, 0) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (380, 0) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (380, 0) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (380, 0) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (380, 0) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (380, 0) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (380, 0) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (380, 0) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (380, 0) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (380, 0) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (380, 0) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (380, 0) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (380, 0) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (380, 0) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (380, 0) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (380, 0) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (380, 0) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (380, 0) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (380, 0) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (380, 0) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (380, 0) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 20
		if (frame_counter == 7'd20 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (400, 0) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (400, 0) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (400, 0) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (400, 0) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (400, 0) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (400, 0) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (400, 0) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (400, 0) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (400, 0) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (400, 0) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (400, 0) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (400, 0) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (400, 0) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (400, 0) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (400, 0) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (400, 0) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (400, 0) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (400, 0) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (400, 0) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (400, 0) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (400, 0) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (400, 0) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (400, 0) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (400, 0) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (400, 0) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (400, 0) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (400, 0) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (400, 0) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (400, 0) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (400, 0) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (400, 0) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (400, 0) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (400, 0) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (400, 0) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (400, 0) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (400, 0) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (400, 0) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (400, 0) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (400, 0) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (400, 0) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (400, 0) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (400, 0) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (400, 0) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (400, 0) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (400, 0) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (400, 0) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (400, 0) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (400, 0) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (400, 0) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (400, 0) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (400, 0) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (400, 0) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (400, 0) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (400, 0) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (400, 0) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (400, 0) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (400, 0) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (400, 0) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (400, 0) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (400, 0) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (400, 0) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (400, 0) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (400, 0) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (400, 0) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (400, 0) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (400, 0) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (400, 0) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (400, 0) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (400, 0) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (400, 0) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (400, 0) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (400, 0) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (400, 0) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (400, 0) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (400, 0) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (400, 0) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (400, 0) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (400, 0) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (400, 0) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (400, 0) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (400, 0) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (400, 0) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (400, 0) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (400, 0) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (400, 0) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (400, 0) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (400, 0) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (400, 0) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (400, 0) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (400, 0) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (400, 0) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (400, 0) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (400, 0) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (400, 0) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (400, 0) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (400, 0) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (400, 0) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (400, 0) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (400, 0) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (400, 0) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (400, 0) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (400, 0) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (400, 0) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (400, 0) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (400, 0) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (400, 0) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (400, 0) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (400, 0) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (400, 0) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (400, 0) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (400, 0) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (400, 0) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 21
		if (frame_counter == 7'd21 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (420, 0) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (420, 0) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (420, 0) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (420, 0) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (420, 0) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (420, 0) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (420, 0) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (420, 0) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (420, 0) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (420, 0) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (420, 0) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (420, 0) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (420, 0) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (420, 0) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (420, 0) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (420, 0) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (420, 0) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (420, 0) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (420, 0) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (420, 0) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (420, 0) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (420, 0) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (420, 0) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (420, 0) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (420, 0) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (420, 0) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (420, 0) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (420, 0) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (420, 0) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (420, 0) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (420, 0) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (420, 0) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (420, 0) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (420, 0) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (420, 0) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (420, 0) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (420, 0) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (420, 0) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (420, 0) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (420, 0) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (420, 0) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (420, 0) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (420, 0) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (420, 0) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (420, 0) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (420, 0) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (420, 0) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (420, 0) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (420, 0) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (420, 0) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (420, 0) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (420, 0) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (420, 0) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (420, 0) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (420, 0) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (420, 0) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (420, 0) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (420, 0) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (420, 0) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (420, 0) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (420, 0) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (420, 0) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (420, 0) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (420, 0) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (420, 0) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (420, 0) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (420, 0) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (420, 0) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (420, 0) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (420, 0) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (420, 0) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (420, 0) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (420, 0) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (420, 0) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (420, 0) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (420, 0) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (420, 0) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (420, 0) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (420, 0) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (420, 0) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (420, 0) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (420, 0) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (420, 0) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (420, 0) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (420, 0) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (420, 0) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (420, 0) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (420, 0) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (420, 0) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (420, 0) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (420, 0) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (420, 0) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (420, 0) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (420, 0) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (420, 0) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (420, 0) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (420, 0) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (420, 0) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (420, 0) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (420, 0) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (420, 0) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (420, 0) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (420, 0) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (420, 0) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (420, 0) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (420, 0) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (420, 0) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (420, 0) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (420, 0) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (420, 0) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (420, 0) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (420, 0) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 22
		if (frame_counter == 7'd22 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (440, 0) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (440, 0) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (440, 0) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (440, 0) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (440, 0) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (440, 0) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (440, 0) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (440, 0) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (440, 0) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (440, 0) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (440, 0) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (440, 0) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (440, 0) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (440, 0) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (440, 0) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (440, 0) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (440, 0) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (440, 0) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (440, 0) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (440, 0) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (440, 0) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (440, 0) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (440, 0) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (440, 0) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (440, 0) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (440, 0) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (440, 0) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (440, 0) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (440, 0) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (440, 0) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (440, 0) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (440, 0) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (440, 0) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (440, 0) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (440, 0) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (440, 0) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (440, 0) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (440, 0) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (440, 0) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (440, 0) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (440, 0) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (440, 0) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (440, 0) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (440, 0) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (440, 0) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (440, 0) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (440, 0) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (440, 0) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (440, 0) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (440, 0) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (440, 0) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (440, 0) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (440, 0) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (440, 0) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (440, 0) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (440, 0) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (440, 0) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (440, 0) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (440, 0) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (440, 0) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (440, 0) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (440, 0) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (440, 0) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (440, 0) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (440, 0) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (440, 0) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (440, 0) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (440, 0) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (440, 0) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (440, 0) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (440, 0) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (440, 0) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (440, 0) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (440, 0) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (440, 0) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (440, 0) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (440, 0) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (440, 0) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (440, 0) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (440, 0) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (440, 0) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (440, 0) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (440, 0) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (440, 0) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (440, 0) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (440, 0) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (440, 0) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (440, 0) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (440, 0) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (440, 0) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (440, 0) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (440, 0) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (440, 0) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (440, 0) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (440, 0) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (440, 0) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (440, 0) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (440, 0) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (440, 0) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (440, 0) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (440, 0) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (440, 0) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (440, 0) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (440, 0) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (440, 0) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (440, 0) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (440, 0) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (440, 0) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (440, 0) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (440, 0) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (440, 0) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (440, 0) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 23
		if (frame_counter == 7'd23 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (460, 0) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (460, 0) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (460, 0) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (460, 0) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (460, 0) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (460, 0) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (460, 0) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (460, 0) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (460, 0) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (460, 0) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (460, 0) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (460, 0) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (460, 0) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (460, 0) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (460, 0) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (460, 0) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (460, 0) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (460, 0) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (460, 0) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (460, 0) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (460, 0) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (460, 0) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (460, 0) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (460, 0) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (460, 0) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (460, 0) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (460, 0) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (460, 0) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (460, 0) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (460, 0) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (460, 0) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (460, 0) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (460, 0) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (460, 0) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (460, 0) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (460, 0) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (460, 0) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (460, 0) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (460, 0) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (460, 0) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (460, 0) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (460, 0) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (460, 0) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (460, 0) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (460, 0) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (460, 0) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (460, 0) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (460, 0) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (460, 0) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (460, 0) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (460, 0) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (460, 0) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (460, 0) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (460, 0) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (460, 0) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (460, 0) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (460, 0) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (460, 0) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (460, 0) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (460, 0) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (460, 0) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (460, 0) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (460, 0) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (460, 0) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (460, 0) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (460, 0) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (460, 0) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (460, 0) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (460, 0) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (460, 0) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (460, 0) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (460, 0) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (460, 0) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (460, 0) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (460, 0) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (460, 0) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (460, 0) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (460, 0) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (460, 0) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (460, 0) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (460, 0) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (460, 0) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (460, 0) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (460, 0) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (460, 0) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (460, 0) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (460, 0) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (460, 0) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (460, 0) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (460, 0) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (460, 0) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (460, 0) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (460, 0) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (460, 0) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (460, 0) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (460, 0) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (460, 0) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (460, 0) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (460, 0) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (460, 0) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (460, 0) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (460, 0) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (460, 0) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (460, 0) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (460, 0) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (460, 0) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (460, 0) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (460, 0) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (460, 0) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (460, 0) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (460, 0) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (460, 0) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 24
		if (frame_counter == 7'd24 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (480, 0) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (480, 0) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (480, 0) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (480, 0) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (480, 0) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (480, 0) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (480, 0) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (480, 0) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (480, 0) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (480, 0) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (480, 0) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (480, 0) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (480, 0) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (480, 0) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (480, 0) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (480, 0) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (480, 0) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (480, 0) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (480, 0) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (480, 0) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (480, 0) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (480, 0) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (480, 0) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (480, 0) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (480, 0) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (480, 0) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (480, 0) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (480, 0) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (480, 0) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (480, 0) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (480, 0) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (480, 0) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (480, 0) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (480, 0) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (480, 0) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (480, 0) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (480, 0) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (480, 0) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (480, 0) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (480, 0) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (480, 0) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (480, 0) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (480, 0) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (480, 0) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (480, 0) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (480, 0) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (480, 0) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (480, 0) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (480, 0) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (480, 0) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (480, 0) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (480, 0) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (480, 0) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (480, 0) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (480, 0) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (480, 0) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (480, 0) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (480, 0) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (480, 0) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (480, 0) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (480, 0) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (480, 0) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (480, 0) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (480, 0) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (480, 0) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (480, 0) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (480, 0) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (480, 0) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (480, 0) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (480, 0) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (480, 0) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (480, 0) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (480, 0) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (480, 0) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (480, 0) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (480, 0) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (480, 0) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (480, 0) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (480, 0) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (480, 0) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (480, 0) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (480, 0) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (480, 0) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (480, 0) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (480, 0) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (480, 0) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (480, 0) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (480, 0) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (480, 0) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (480, 0) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (480, 0) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (480, 0) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (480, 0) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (480, 0) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (480, 0) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (480, 0) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (480, 0) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (480, 0) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (480, 0) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (480, 0) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (480, 0) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (480, 0) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (480, 0) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (480, 0) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (480, 0) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (480, 0) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (480, 0) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (480, 0) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (480, 0) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (480, 0) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (480, 0) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (480, 0) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 25
		if (frame_counter == 7'd25 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (500, 0) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (500, 0) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (500, 0) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (500, 0) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (500, 0) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (500, 0) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (500, 0) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (500, 0) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (500, 0) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (500, 0) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (500, 0) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (500, 0) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (500, 0) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (500, 0) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (500, 0) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (500, 0) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (500, 0) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (500, 0) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (500, 0) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (500, 0) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (500, 0) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (500, 0) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (500, 0) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (500, 0) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (500, 0) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (500, 0) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (500, 0) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (500, 0) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (500, 0) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (500, 0) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (500, 0) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (500, 0) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (500, 0) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (500, 0) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (500, 0) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (500, 0) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (500, 0) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (500, 0) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (500, 0) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (500, 0) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (500, 0) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (500, 0) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (500, 0) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (500, 0) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (500, 0) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (500, 0) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (500, 0) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (500, 0) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (500, 0) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (500, 0) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (500, 0) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (500, 0) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (500, 0) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (500, 0) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (500, 0) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (500, 0) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (500, 0) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (500, 0) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (500, 0) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (500, 0) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (500, 0) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (500, 0) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (500, 0) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (500, 0) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (500, 0) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (500, 0) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (500, 0) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (500, 0) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (500, 0) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (500, 0) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (500, 0) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (500, 0) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (500, 0) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (500, 0) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (500, 0) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (500, 0) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (500, 0) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (500, 0) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (500, 0) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (500, 0) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (500, 0) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (500, 0) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (500, 0) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (500, 0) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (500, 0) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (500, 0) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (500, 0) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (500, 0) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (500, 0) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (500, 0) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (500, 0) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (500, 0) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (500, 0) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (500, 0) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (500, 0) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (500, 0) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (500, 0) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (500, 0) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (500, 0) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (500, 0) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (500, 0) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (500, 0) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (500, 0) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (500, 0) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (500, 0) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (500, 0) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (500, 0) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (500, 0) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (500, 0) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (500, 0) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (500, 0) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (500, 0) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 26
		if (frame_counter == 7'd26 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (520, 0) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (520, 0) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (520, 0) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (520, 0) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (520, 0) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (520, 0) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (520, 0) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (520, 0) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (520, 0) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (520, 0) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (520, 0) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (520, 0) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (520, 0) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (520, 0) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (520, 0) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (520, 0) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (520, 0) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (520, 0) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (520, 0) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (520, 0) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (520, 0) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (520, 0) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (520, 0) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (520, 0) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (520, 0) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (520, 0) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (520, 0) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (520, 0) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (520, 0) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (520, 0) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (520, 0) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (520, 0) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (520, 0) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (520, 0) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (520, 0) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (520, 0) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (520, 0) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (520, 0) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (520, 0) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (520, 0) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (520, 0) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (520, 0) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (520, 0) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (520, 0) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (520, 0) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (520, 0) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (520, 0) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (520, 0) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (520, 0) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (520, 0) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (520, 0) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (520, 0) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (520, 0) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (520, 0) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (520, 0) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (520, 0) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (520, 0) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (520, 0) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (520, 0) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (520, 0) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (520, 0) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (520, 0) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (520, 0) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (520, 0) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (520, 0) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (520, 0) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (520, 0) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (520, 0) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (520, 0) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (520, 0) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (520, 0) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (520, 0) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (520, 0) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (520, 0) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (520, 0) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (520, 0) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (520, 0) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (520, 0) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (520, 0) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (520, 0) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (520, 0) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (520, 0) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (520, 0) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (520, 0) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (520, 0) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (520, 0) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (520, 0) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (520, 0) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (520, 0) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (520, 0) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (520, 0) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (520, 0) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (520, 0) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (520, 0) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (520, 0) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (520, 0) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (520, 0) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (520, 0) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (520, 0) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (520, 0) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (520, 0) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (520, 0) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (520, 0) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (520, 0) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (520, 0) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (520, 0) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (520, 0) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (520, 0) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (520, 0) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (520, 0) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (520, 0) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (520, 0) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 27
		if (frame_counter == 7'd27 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (540, 0) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (540, 0) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (540, 0) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (540, 0) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (540, 0) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (540, 0) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (540, 0) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (540, 0) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (540, 0) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (540, 0) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (540, 0) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (540, 0) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (540, 0) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (540, 0) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (540, 0) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (540, 0) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (540, 0) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (540, 0) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (540, 0) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (540, 0) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (540, 0) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (540, 0) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (540, 0) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (540, 0) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (540, 0) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (540, 0) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (540, 0) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (540, 0) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (540, 0) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (540, 0) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (540, 0) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (540, 0) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (540, 0) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (540, 0) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (540, 0) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (540, 0) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (540, 0) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (540, 0) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (540, 0) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (540, 0) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (540, 0) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (540, 0) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (540, 0) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (540, 0) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (540, 0) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (540, 0) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (540, 0) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (540, 0) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (540, 0) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (540, 0) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (540, 0) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (540, 0) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (540, 0) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (540, 0) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (540, 0) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (540, 0) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (540, 0) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (540, 0) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (540, 0) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (540, 0) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (540, 0) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (540, 0) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (540, 0) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (540, 0) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (540, 0) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (540, 0) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (540, 0) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (540, 0) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (540, 0) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (540, 0) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (540, 0) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (540, 0) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (540, 0) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (540, 0) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (540, 0) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (540, 0) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (540, 0) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (540, 0) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (540, 0) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (540, 0) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (540, 0) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (540, 0) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (540, 0) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (540, 0) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (540, 0) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (540, 0) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (540, 0) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (540, 0) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (540, 0) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (540, 0) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (540, 0) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (540, 0) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (540, 0) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (540, 0) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (540, 0) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (540, 0) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (540, 0) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (540, 0) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (540, 0) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (540, 0) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (540, 0) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (540, 0) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (540, 0) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (540, 0) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (540, 0) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (540, 0) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (540, 0) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (540, 0) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (540, 0) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (540, 0) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (540, 0) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (540, 0) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 28
		if (frame_counter == 7'd28 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (560, 0) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (560, 0) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (560, 0) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (560, 0) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (560, 0) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (560, 0) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (560, 0) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (560, 0) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (560, 0) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (560, 0) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (560, 0) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (560, 0) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (560, 0) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (560, 0) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (560, 0) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (560, 0) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (560, 0) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (560, 0) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (560, 0) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (560, 0) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (560, 0) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (560, 0) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (560, 0) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (560, 0) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (560, 0) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (560, 0) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (560, 0) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (560, 0) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (560, 0) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (560, 0) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (560, 0) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (560, 0) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (560, 0) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (560, 0) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (560, 0) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (560, 0) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (560, 0) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (560, 0) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (560, 0) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (560, 0) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (560, 0) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (560, 0) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (560, 0) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (560, 0) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (560, 0) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (560, 0) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (560, 0) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (560, 0) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (560, 0) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (560, 0) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (560, 0) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (560, 0) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (560, 0) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (560, 0) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (560, 0) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (560, 0) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (560, 0) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (560, 0) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (560, 0) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (560, 0) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (560, 0) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (560, 0) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (560, 0) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (560, 0) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (560, 0) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (560, 0) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (560, 0) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (560, 0) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (560, 0) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (560, 0) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (560, 0) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (560, 0) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (560, 0) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (560, 0) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (560, 0) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (560, 0) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (560, 0) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (560, 0) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (560, 0) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (560, 0) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (560, 0) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (560, 0) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (560, 0) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (560, 0) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (560, 0) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (560, 0) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (560, 0) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (560, 0) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (560, 0) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (560, 0) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (560, 0) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (560, 0) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (560, 0) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (560, 0) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (560, 0) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (560, 0) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (560, 0) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (560, 0) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (560, 0) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (560, 0) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (560, 0) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (560, 0) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (560, 0) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (560, 0) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (560, 0) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (560, 0) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (560, 0) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (560, 0) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (560, 0) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (560, 0) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (560, 0) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (560, 0) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 29
		if (frame_counter == 7'd29 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (580, 0) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (580, 0) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (580, 0) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (580, 0) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (580, 0) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (580, 0) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (580, 0) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (580, 0) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (580, 0) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (580, 0) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (580, 0) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (580, 0) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (580, 0) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (580, 0) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (580, 0) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (580, 0) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (580, 0) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (580, 0) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (580, 0) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (580, 0) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (580, 0) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (580, 0) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (580, 0) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (580, 0) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (580, 0) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (580, 0) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (580, 0) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (580, 0) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (580, 0) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (580, 0) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (580, 0) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (580, 0) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (580, 0) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (580, 0) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (580, 0) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (580, 0) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (580, 0) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (580, 0) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (580, 0) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (580, 0) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (580, 0) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (580, 0) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (580, 0) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (580, 0) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (580, 0) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (580, 0) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (580, 0) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (580, 0) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (580, 0) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (580, 0) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (580, 0) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (580, 0) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (580, 0) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (580, 0) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (580, 0) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (580, 0) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (580, 0) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (580, 0) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (580, 0) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (580, 0) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (580, 0) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (580, 0) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (580, 0) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (580, 0) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (580, 0) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (580, 0) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (580, 0) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (580, 0) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (580, 0) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (580, 0) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (580, 0) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (580, 0) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (580, 0) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (580, 0) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (580, 0) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (580, 0) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (580, 0) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (580, 0) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (580, 0) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (580, 0) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (580, 0) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (580, 0) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (580, 0) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (580, 0) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (580, 0) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (580, 0) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (580, 0) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (580, 0) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (580, 0) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (580, 0) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (580, 0) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (580, 0) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (580, 0) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (580, 0) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (580, 0) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (580, 0) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (580, 0) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (580, 0) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (580, 0) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (580, 0) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (580, 0) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (580, 0) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (580, 0) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (580, 0) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (580, 0) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (580, 0) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (580, 0) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (580, 0) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (580, 0) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (580, 0) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (580, 0) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (580, 0) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 30
		if (frame_counter == 7'd30 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (600, 0) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (600, 0) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (600, 0) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (600, 0) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (600, 0) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (600, 0) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (600, 0) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (600, 0) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (600, 0) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (600, 0) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (600, 0) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (600, 0) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (600, 0) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (600, 0) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (600, 0) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (600, 0) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (600, 0) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (600, 0) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (600, 0) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (600, 0) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (600, 0) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (600, 0) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (600, 0) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (600, 0) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (600, 0) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (600, 0) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (600, 0) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (600, 0) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (600, 0) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (600, 0) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (600, 0) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (600, 0) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (600, 0) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (600, 0) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (600, 0) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (600, 0) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (600, 0) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (600, 0) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (600, 0) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (600, 0) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (600, 0) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (600, 0) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (600, 0) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (600, 0) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (600, 0) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (600, 0) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (600, 0) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (600, 0) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (600, 0) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (600, 0) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (600, 0) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (600, 0) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (600, 0) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (600, 0) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (600, 0) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (600, 0) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (600, 0) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (600, 0) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (600, 0) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (600, 0) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (600, 0) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (600, 0) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (600, 0) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (600, 0) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (600, 0) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (600, 0) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (600, 0) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (600, 0) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (600, 0) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (600, 0) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (600, 0) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (600, 0) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (600, 0) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (600, 0) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (600, 0) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (600, 0) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (600, 0) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (600, 0) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (600, 0) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (600, 0) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (600, 0) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (600, 0) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (600, 0) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (600, 0) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (600, 0) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (600, 0) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (600, 0) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (600, 0) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (600, 0) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (600, 0) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (600, 0) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (600, 0) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (600, 0) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (600, 0) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (600, 0) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (600, 0) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (600, 0) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (600, 0) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (600, 0) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (600, 0) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (600, 0) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (600, 0) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (600, 0) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (600, 0) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (600, 0) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (600, 0) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (600, 0) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (600, 0) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (600, 0) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (600, 0) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (600, 0) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (600, 0) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 31
		if (frame_counter == 7'd31 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (620, 0) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (620, 0) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (620, 0) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (620, 0) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (620, 0) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (620, 0) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (620, 0) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (620, 0) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (620, 0) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (620, 0) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (620, 0) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (620, 0) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (620, 0) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (620, 0) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (620, 0) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (620, 0) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (620, 0) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (620, 0) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (620, 0) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (620, 0) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (620, 0) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (620, 0) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (620, 0) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (620, 0) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (620, 0) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (620, 0) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (620, 0) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (620, 0) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (620, 0) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (620, 0) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (620, 0) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (620, 0) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (620, 0) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (620, 0) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (620, 0) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (620, 0) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (620, 0) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (620, 0) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (620, 0) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (620, 0) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (620, 0) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (620, 0) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (620, 0) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (620, 0) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (620, 0) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (620, 0) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (620, 0) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (620, 0) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (620, 0) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (620, 0) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (620, 0) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (620, 0) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (620, 0) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (620, 0) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (620, 0) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (620, 0) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (620, 0) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (620, 0) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (620, 0) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (620, 0) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (620, 0) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (620, 0) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (620, 0) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (620, 0) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (620, 0) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (620, 0) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (620, 0) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (620, 0) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (620, 0) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (620, 0) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (620, 0) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (620, 0) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (620, 0) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (620, 0) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (620, 0) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (620, 0) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (620, 0) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (620, 0) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (620, 0) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (620, 0) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (620, 0) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (620, 0) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (620, 0) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (620, 0) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (620, 0) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (620, 0) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (620, 0) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (620, 0) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (620, 0) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (620, 0) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (620, 0) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (620, 0) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (620, 0) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (620, 0) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (620, 0) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (620, 0) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (620, 0) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (620, 0) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (620, 0) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (620, 0) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (620, 0) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (620, 0) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (620, 0) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (620, 0) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (620, 0) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (620, 0) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (620, 0) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (620, 0) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (620, 0) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (620, 0) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (620, 0) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (620, 0) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 32
		if (frame_counter == 7'd32 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (640, 0) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (640, 0) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (640, 0) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (640, 0) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (640, 0) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (640, 0) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (640, 0) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (640, 0) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (640, 0) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (640, 0) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (640, 0) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (640, 0) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (640, 0) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (640, 0) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (640, 0) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (640, 0) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (640, 0) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (640, 0) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (640, 0) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (640, 0) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (640, 0) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (640, 0) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (640, 0) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (640, 0) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (640, 0) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (640, 0) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (640, 0) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (640, 0) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (640, 0) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (640, 0) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (640, 0) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (640, 0) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (640, 0) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (640, 0) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (640, 0) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (640, 0) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (640, 0) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (640, 0) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (640, 0) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (640, 0) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (640, 0) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (640, 0) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (640, 0) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (640, 0) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (640, 0) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (640, 0) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (640, 0) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (640, 0) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (640, 0) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (640, 0) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (640, 0) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (640, 0) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (640, 0) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (640, 0) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (640, 0) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (640, 0) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (640, 0) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (640, 0) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (640, 0) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (640, 0) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (640, 0) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (640, 0) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (640, 0) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (640, 0) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (640, 0) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (640, 0) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (640, 0) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (640, 0) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (640, 0) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (640, 0) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (640, 0) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (640, 0) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (640, 0) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (640, 0) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (640, 0) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (640, 0) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (640, 0) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (640, 0) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (640, 0) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (640, 0) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (640, 0) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (640, 0) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (640, 0) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (640, 0) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (640, 0) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (640, 0) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (640, 0) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (640, 0) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (640, 0) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (640, 0) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (640, 0) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (640, 0) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (640, 0) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (640, 0) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (640, 0) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (640, 0) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (640, 0) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (640, 0) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (640, 0) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (640, 0) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (640, 0) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (640, 0) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (640, 0) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (640, 0) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (640, 0) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (640, 0) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (640, 0) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (640, 0) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (640, 0) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (640, 0) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (640, 0) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (640, 0) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd0;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 33
		if (frame_counter == 7'd33 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (640, 20) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (640, 20) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (640, 20) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (640, 20) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (640, 20) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (640, 20) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (640, 20) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (640, 20) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (640, 20) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (640, 20) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (640, 20) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (640, 20) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (640, 20) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (640, 20) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (640, 20) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (640, 20) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (640, 20) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (640, 20) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (640, 20) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (640, 20) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (640, 20) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (640, 20) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (640, 20) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (640, 20) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (640, 20) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (640, 20) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (640, 20) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (640, 20) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (640, 20) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (640, 20) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (640, 20) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (640, 20) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (640, 20) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (640, 20) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (640, 20) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (640, 20) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (640, 20) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (640, 20) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (640, 20) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (640, 20) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (640, 20) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (640, 20) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (640, 20) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (640, 20) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (640, 20) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (640, 20) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (640, 20) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (640, 20) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (640, 20) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (640, 20) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (640, 20) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (640, 20) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (640, 20) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (640, 20) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (640, 20) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (640, 20) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (640, 20) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (640, 20) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (640, 20) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (640, 20) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (640, 20) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (640, 20) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (640, 20) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (640, 20) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (640, 20) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (640, 20) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (640, 20) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (640, 20) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (640, 20) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (640, 20) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (640, 20) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (640, 20) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (640, 20) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (640, 20) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (640, 20) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (640, 20) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (640, 20) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (640, 20) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (640, 20) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (640, 20) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (640, 20) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (640, 20) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (640, 20) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (640, 20) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (640, 20) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (640, 20) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (640, 20) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (640, 20) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (640, 20) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (640, 20) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (640, 20) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (640, 20) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (640, 20) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (640, 20) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (640, 20) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (640, 20) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (640, 20) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (640, 20) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (640, 20) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (640, 20) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (640, 20) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (640, 20) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (640, 20) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (640, 20) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (640, 20) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (640, 20) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (640, 20) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (640, 20) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (640, 20) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (640, 20) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (640, 20) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (640, 20) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd20;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 34
		if (frame_counter == 7'd34 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (640, 40) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (640, 40) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (640, 40) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (640, 40) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (640, 40) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (640, 40) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (640, 40) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (640, 40) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (640, 40) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (640, 40) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (640, 40) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (640, 40) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (640, 40) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (640, 40) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (640, 40) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (640, 40) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (640, 40) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (640, 40) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (640, 40) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (640, 40) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (640, 40) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (640, 40) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (640, 40) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (640, 40) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (640, 40) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (640, 40) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (640, 40) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (640, 40) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (640, 40) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (640, 40) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (640, 40) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (640, 40) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (640, 40) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (640, 40) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (640, 40) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (640, 40) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (640, 40) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (640, 40) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (640, 40) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (640, 40) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (640, 40) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (640, 40) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (640, 40) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (640, 40) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (640, 40) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (640, 40) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (640, 40) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (640, 40) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (640, 40) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (640, 40) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (640, 40) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (640, 40) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (640, 40) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (640, 40) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (640, 40) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (640, 40) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (640, 40) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (640, 40) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (640, 40) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (640, 40) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (640, 40) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (640, 40) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (640, 40) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (640, 40) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (640, 40) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (640, 40) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (640, 40) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (640, 40) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (640, 40) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (640, 40) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (640, 40) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (640, 40) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (640, 40) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (640, 40) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (640, 40) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (640, 40) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (640, 40) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (640, 40) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (640, 40) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (640, 40) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (640, 40) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (640, 40) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (640, 40) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (640, 40) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (640, 40) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (640, 40) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (640, 40) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (640, 40) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (640, 40) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (640, 40) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (640, 40) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (640, 40) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (640, 40) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (640, 40) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (640, 40) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (640, 40) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (640, 40) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (640, 40) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (640, 40) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (640, 40) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (640, 40) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (640, 40) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (640, 40) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (640, 40) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (640, 40) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (640, 40) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (640, 40) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (640, 40) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (640, 40) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (640, 40) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (640, 40) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (640, 40) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd40;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 35
		if (frame_counter == 7'd35 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (640, 60) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (640, 60) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (640, 60) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (640, 60) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (640, 60) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (640, 60) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (640, 60) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (640, 60) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (640, 60) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (640, 60) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (640, 60) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (640, 60) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (640, 60) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (640, 60) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (640, 60) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (640, 60) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (640, 60) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (640, 60) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (640, 60) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (640, 60) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (640, 60) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (640, 60) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (640, 60) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (640, 60) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (640, 60) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (640, 60) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (640, 60) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (640, 60) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (640, 60) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (640, 60) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (640, 60) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (640, 60) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (640, 60) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (640, 60) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (640, 60) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (640, 60) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (640, 60) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (640, 60) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (640, 60) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (640, 60) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (640, 60) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (640, 60) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (640, 60) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (640, 60) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (640, 60) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (640, 60) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (640, 60) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (640, 60) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (640, 60) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (640, 60) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (640, 60) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (640, 60) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (640, 60) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (640, 60) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (640, 60) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (640, 60) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (640, 60) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (640, 60) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (640, 60) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (640, 60) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (640, 60) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (640, 60) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (640, 60) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (640, 60) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (640, 60) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (640, 60) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (640, 60) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (640, 60) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (640, 60) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (640, 60) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (640, 60) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (640, 60) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (640, 60) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (640, 60) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (640, 60) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (640, 60) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (640, 60) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (640, 60) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (640, 60) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (640, 60) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (640, 60) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (640, 60) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (640, 60) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (640, 60) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (640, 60) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (640, 60) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (640, 60) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (640, 60) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (640, 60) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (640, 60) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (640, 60) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (640, 60) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (640, 60) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (640, 60) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (640, 60) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (640, 60) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (640, 60) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (640, 60) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (640, 60) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (640, 60) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (640, 60) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (640, 60) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (640, 60) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (640, 60) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (640, 60) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (640, 60) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (640, 60) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (640, 60) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (640, 60) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (640, 60) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (640, 60) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (640, 60) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd60;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 36
		if (frame_counter == 7'd36 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (640, 80) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (640, 80) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (640, 80) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (640, 80) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (640, 80) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (640, 80) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (640, 80) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (640, 80) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (640, 80) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (640, 80) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (640, 80) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (640, 80) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (640, 80) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (640, 80) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (640, 80) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (640, 80) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (640, 80) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (640, 80) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (640, 80) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (640, 80) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (640, 80) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (640, 80) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (640, 80) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (640, 80) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (640, 80) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (640, 80) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (640, 80) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (640, 80) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (640, 80) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (640, 80) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (640, 80) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (640, 80) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (640, 80) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (640, 80) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (640, 80) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (640, 80) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (640, 80) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (640, 80) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (640, 80) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (640, 80) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (640, 80) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (640, 80) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (640, 80) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (640, 80) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (640, 80) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (640, 80) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (640, 80) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (640, 80) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (640, 80) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (640, 80) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (640, 80) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (640, 80) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (640, 80) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (640, 80) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (640, 80) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (640, 80) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (640, 80) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (640, 80) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (640, 80) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (640, 80) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (640, 80) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (640, 80) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (640, 80) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (640, 80) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (640, 80) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (640, 80) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (640, 80) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (640, 80) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (640, 80) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (640, 80) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (640, 80) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (640, 80) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (640, 80) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (640, 80) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (640, 80) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (640, 80) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (640, 80) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (640, 80) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (640, 80) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (640, 80) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (640, 80) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (640, 80) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (640, 80) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (640, 80) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (640, 80) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (640, 80) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (640, 80) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (640, 80) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (640, 80) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (640, 80) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (640, 80) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (640, 80) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (640, 80) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (640, 80) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (640, 80) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (640, 80) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (640, 80) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (640, 80) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (640, 80) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (640, 80) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (640, 80) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (640, 80) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (640, 80) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (640, 80) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (640, 80) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (640, 80) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (640, 80) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (640, 80) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (640, 80) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (640, 80) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (640, 80) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (640, 80) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd80;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 37
		if (frame_counter == 7'd37 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (640, 100) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (640, 100) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (640, 100) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (640, 100) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (640, 100) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (640, 100) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (640, 100) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (640, 100) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (640, 100) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (640, 100) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (640, 100) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (640, 100) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (640, 100) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (640, 100) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (640, 100) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (640, 100) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (640, 100) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (640, 100) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (640, 100) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (640, 100) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (640, 100) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (640, 100) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (640, 100) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (640, 100) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (640, 100) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (640, 100) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (640, 100) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (640, 100) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (640, 100) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (640, 100) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (640, 100) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (640, 100) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (640, 100) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (640, 100) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (640, 100) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (640, 100) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (640, 100) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (640, 100) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (640, 100) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (640, 100) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (640, 100) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (640, 100) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (640, 100) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (640, 100) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (640, 100) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (640, 100) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (640, 100) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (640, 100) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (640, 100) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (640, 100) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (640, 100) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (640, 100) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (640, 100) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (640, 100) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (640, 100) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (640, 100) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (640, 100) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (640, 100) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (640, 100) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (640, 100) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (640, 100) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (640, 100) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (640, 100) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (640, 100) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (640, 100) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (640, 100) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (640, 100) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (640, 100) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (640, 100) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (640, 100) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (640, 100) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (640, 100) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (640, 100) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (640, 100) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (640, 100) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (640, 100) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (640, 100) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (640, 100) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (640, 100) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (640, 100) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (640, 100) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (640, 100) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (640, 100) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (640, 100) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (640, 100) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (640, 100) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (640, 100) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (640, 100) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (640, 100) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (640, 100) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (640, 100) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (640, 100) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (640, 100) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (640, 100) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (640, 100) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (640, 100) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (640, 100) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (640, 100) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (640, 100) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (640, 100) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (640, 100) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (640, 100) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (640, 100) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (640, 100) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (640, 100) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (640, 100) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (640, 100) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (640, 100) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (640, 100) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (640, 100) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (640, 100) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (640, 100) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd100;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 38
		if (frame_counter == 7'd38 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (640, 120) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (640, 120) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (640, 120) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (640, 120) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (640, 120) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (640, 120) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (640, 120) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (640, 120) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (640, 120) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (640, 120) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (640, 120) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (640, 120) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (640, 120) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (640, 120) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (640, 120) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (640, 120) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (640, 120) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (640, 120) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (640, 120) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (640, 120) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (640, 120) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (640, 120) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (640, 120) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (640, 120) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (640, 120) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (640, 120) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (640, 120) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (640, 120) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (640, 120) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (640, 120) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (640, 120) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (640, 120) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (640, 120) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (640, 120) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (640, 120) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (640, 120) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (640, 120) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (640, 120) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (640, 120) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (640, 120) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (640, 120) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (640, 120) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (640, 120) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (640, 120) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (640, 120) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (640, 120) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (640, 120) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (640, 120) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (640, 120) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (640, 120) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (640, 120) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (640, 120) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (640, 120) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (640, 120) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (640, 120) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (640, 120) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (640, 120) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (640, 120) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (640, 120) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (640, 120) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (640, 120) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (640, 120) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (640, 120) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (640, 120) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (640, 120) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (640, 120) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (640, 120) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (640, 120) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (640, 120) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (640, 120) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (640, 120) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (640, 120) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (640, 120) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (640, 120) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (640, 120) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (640, 120) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (640, 120) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (640, 120) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (640, 120) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (640, 120) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (640, 120) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (640, 120) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (640, 120) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (640, 120) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (640, 120) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (640, 120) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (640, 120) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (640, 120) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (640, 120) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (640, 120) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (640, 120) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (640, 120) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (640, 120) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (640, 120) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (640, 120) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (640, 120) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (640, 120) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (640, 120) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (640, 120) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (640, 120) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (640, 120) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (640, 120) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (640, 120) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (640, 120) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (640, 120) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (640, 120) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (640, 120) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (640, 120) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (640, 120) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (640, 120) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (640, 120) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (640, 120) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd120;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 39
		if (frame_counter == 7'd39 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (640, 140) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (640, 140) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (640, 140) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (640, 140) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (640, 140) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (640, 140) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (640, 140) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (640, 140) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (640, 140) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (640, 140) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (640, 140) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (640, 140) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (640, 140) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (640, 140) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (640, 140) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (640, 140) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (640, 140) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (640, 140) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (640, 140) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (640, 140) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (640, 140) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (640, 140) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (640, 140) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (640, 140) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (640, 140) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (640, 140) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (640, 140) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (640, 140) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (640, 140) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (640, 140) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (640, 140) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (640, 140) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (640, 140) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (640, 140) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (640, 140) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (640, 140) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (640, 140) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (640, 140) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (640, 140) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (640, 140) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (640, 140) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (640, 140) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (640, 140) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (640, 140) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (640, 140) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (640, 140) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (640, 140) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (640, 140) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (640, 140) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (640, 140) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (640, 140) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (640, 140) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (640, 140) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (640, 140) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (640, 140) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (640, 140) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (640, 140) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (640, 140) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (640, 140) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (640, 140) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (640, 140) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (640, 140) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (640, 140) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (640, 140) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (640, 140) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (640, 140) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (640, 140) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (640, 140) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (640, 140) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (640, 140) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (640, 140) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (640, 140) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (640, 140) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (640, 140) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (640, 140) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (640, 140) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (640, 140) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (640, 140) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (640, 140) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (640, 140) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (640, 140) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (640, 140) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (640, 140) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (640, 140) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (640, 140) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (640, 140) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (640, 140) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (640, 140) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (640, 140) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (640, 140) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (640, 140) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (640, 140) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (640, 140) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (640, 140) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (640, 140) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (640, 140) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (640, 140) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (640, 140) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (640, 140) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (640, 140) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (640, 140) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (640, 140) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (640, 140) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (640, 140) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (640, 140) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (640, 140) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (640, 140) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (640, 140) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (640, 140) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (640, 140) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (640, 140) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (640, 140) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd140;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 40
		if (frame_counter == 7'd40 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (640, 160) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (640, 160) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (640, 160) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (640, 160) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (640, 160) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (640, 160) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (640, 160) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (640, 160) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (640, 160) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (640, 160) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (640, 160) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (640, 160) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (640, 160) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (640, 160) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (640, 160) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (640, 160) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (640, 160) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (640, 160) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (640, 160) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (640, 160) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (640, 160) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (640, 160) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (640, 160) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (640, 160) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (640, 160) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (640, 160) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (640, 160) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (640, 160) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (640, 160) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (640, 160) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (640, 160) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (640, 160) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (640, 160) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (640, 160) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (640, 160) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (640, 160) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (640, 160) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (640, 160) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (640, 160) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (640, 160) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (640, 160) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (640, 160) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (640, 160) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (640, 160) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (640, 160) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (640, 160) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (640, 160) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (640, 160) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (640, 160) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (640, 160) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (640, 160) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (640, 160) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (640, 160) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (640, 160) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (640, 160) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (640, 160) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (640, 160) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (640, 160) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (640, 160) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (640, 160) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (640, 160) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (640, 160) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (640, 160) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (640, 160) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (640, 160) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (640, 160) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (640, 160) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (640, 160) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (640, 160) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (640, 160) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (640, 160) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (640, 160) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (640, 160) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (640, 160) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (640, 160) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (640, 160) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (640, 160) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (640, 160) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (640, 160) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (640, 160) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (640, 160) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (640, 160) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (640, 160) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (640, 160) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (640, 160) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (640, 160) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (640, 160) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (640, 160) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (640, 160) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (640, 160) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (640, 160) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (640, 160) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (640, 160) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (640, 160) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (640, 160) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (640, 160) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (640, 160) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (640, 160) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (640, 160) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (640, 160) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (640, 160) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (640, 160) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (640, 160) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (640, 160) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (640, 160) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (640, 160) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (640, 160) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (640, 160) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (640, 160) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (640, 160) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (640, 160) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (640, 160) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd160;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 41
		if (frame_counter == 7'd41 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (640, 180) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (640, 180) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (640, 180) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (640, 180) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (640, 180) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (640, 180) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (640, 180) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (640, 180) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (640, 180) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (640, 180) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (640, 180) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (640, 180) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (640, 180) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (640, 180) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (640, 180) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (640, 180) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (640, 180) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (640, 180) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (640, 180) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (640, 180) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (640, 180) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (640, 180) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (640, 180) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (640, 180) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (640, 180) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (640, 180) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (640, 180) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (640, 180) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (640, 180) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (640, 180) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (640, 180) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (640, 180) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (640, 180) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (640, 180) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (640, 180) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (640, 180) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (640, 180) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (640, 180) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (640, 180) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (640, 180) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (640, 180) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (640, 180) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (640, 180) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (640, 180) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (640, 180) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (640, 180) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (640, 180) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (640, 180) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (640, 180) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (640, 180) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (640, 180) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (640, 180) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (640, 180) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (640, 180) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (640, 180) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (640, 180) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (640, 180) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (640, 180) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (640, 180) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (640, 180) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (640, 180) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (640, 180) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (640, 180) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (640, 180) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (640, 180) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (640, 180) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (640, 180) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (640, 180) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (640, 180) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (640, 180) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (640, 180) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (640, 180) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (640, 180) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (640, 180) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (640, 180) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (640, 180) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (640, 180) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (640, 180) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (640, 180) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (640, 180) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (640, 180) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (640, 180) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (640, 180) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (640, 180) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (640, 180) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (640, 180) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (640, 180) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (640, 180) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (640, 180) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (640, 180) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (640, 180) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (640, 180) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (640, 180) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (640, 180) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (640, 180) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (640, 180) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (640, 180) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (640, 180) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (640, 180) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (640, 180) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (640, 180) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (640, 180) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (640, 180) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (640, 180) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (640, 180) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (640, 180) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (640, 180) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (640, 180) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (640, 180) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (640, 180) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (640, 180) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (640, 180) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd180;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 42
		if (frame_counter == 7'd42 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (640, 200) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (640, 200) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (640, 200) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (640, 200) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (640, 200) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (640, 200) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (640, 200) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (640, 200) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (640, 200) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (640, 200) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (640, 200) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (640, 200) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (640, 200) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (640, 200) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (640, 200) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (640, 200) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (640, 200) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (640, 200) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (640, 200) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (640, 200) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (640, 200) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (640, 200) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (640, 200) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (640, 200) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (640, 200) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (640, 200) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (640, 200) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (640, 200) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (640, 200) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (640, 200) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (640, 200) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (640, 200) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (640, 200) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (640, 200) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (640, 200) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (640, 200) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (640, 200) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (640, 200) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (640, 200) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (640, 200) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (640, 200) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (640, 200) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (640, 200) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (640, 200) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (640, 200) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (640, 200) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (640, 200) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (640, 200) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (640, 200) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (640, 200) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (640, 200) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (640, 200) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (640, 200) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (640, 200) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (640, 200) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (640, 200) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (640, 200) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (640, 200) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (640, 200) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (640, 200) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (640, 200) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (640, 200) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (640, 200) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (640, 200) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (640, 200) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (640, 200) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (640, 200) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (640, 200) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (640, 200) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (640, 200) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (640, 200) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (640, 200) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (640, 200) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (640, 200) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (640, 200) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (640, 200) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (640, 200) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (640, 200) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (640, 200) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (640, 200) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (640, 200) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (640, 200) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (640, 200) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (640, 200) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (640, 200) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (640, 200) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (640, 200) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (640, 200) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (640, 200) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (640, 200) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (640, 200) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (640, 200) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (640, 200) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (640, 200) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (640, 200) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (640, 200) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (640, 200) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (640, 200) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (640, 200) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (640, 200) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (640, 200) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (640, 200) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (640, 200) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (640, 200) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (640, 200) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (640, 200) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (640, 200) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (640, 200) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (640, 200) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (640, 200) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (640, 200) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (640, 200) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd200;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 43
		if (frame_counter == 7'd43 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (640, 220) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (640, 220) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (640, 220) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (640, 220) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (640, 220) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (640, 220) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (640, 220) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (640, 220) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (640, 220) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (640, 220) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (640, 220) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (640, 220) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (640, 220) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (640, 220) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (640, 220) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (640, 220) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (640, 220) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (640, 220) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (640, 220) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (640, 220) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (640, 220) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (640, 220) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (640, 220) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (640, 220) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (640, 220) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (640, 220) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (640, 220) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (640, 220) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (640, 220) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (640, 220) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (640, 220) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (640, 220) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (640, 220) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (640, 220) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (640, 220) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (640, 220) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (640, 220) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (640, 220) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (640, 220) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (640, 220) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (640, 220) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (640, 220) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (640, 220) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (640, 220) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (640, 220) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (640, 220) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (640, 220) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (640, 220) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (640, 220) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (640, 220) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (640, 220) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (640, 220) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (640, 220) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (640, 220) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (640, 220) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (640, 220) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (640, 220) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (640, 220) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (640, 220) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (640, 220) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (640, 220) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (640, 220) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (640, 220) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (640, 220) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (640, 220) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (640, 220) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (640, 220) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (640, 220) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (640, 220) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (640, 220) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (640, 220) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (640, 220) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (640, 220) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (640, 220) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (640, 220) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (640, 220) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (640, 220) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (640, 220) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (640, 220) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (640, 220) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (640, 220) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (640, 220) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (640, 220) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (640, 220) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (640, 220) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (640, 220) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (640, 220) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (640, 220) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (640, 220) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (640, 220) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (640, 220) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (640, 220) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (640, 220) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (640, 220) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (640, 220) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (640, 220) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (640, 220) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (640, 220) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (640, 220) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (640, 220) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (640, 220) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (640, 220) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (640, 220) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (640, 220) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (640, 220) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (640, 220) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (640, 220) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (640, 220) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (640, 220) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (640, 220) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (640, 220) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (640, 220) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd220;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 44
		if (frame_counter == 7'd44 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (640, 240) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (640, 240) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (640, 240) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (640, 240) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (640, 240) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (640, 240) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (640, 240) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (640, 240) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (640, 240) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (640, 240) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (640, 240) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (640, 240) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (640, 240) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (640, 240) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (640, 240) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (640, 240) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (640, 240) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (640, 240) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (640, 240) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (640, 240) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (640, 240) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (640, 240) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (640, 240) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (640, 240) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (640, 240) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (640, 240) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (640, 240) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (640, 240) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (640, 240) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (640, 240) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (640, 240) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (640, 240) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (640, 240) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (640, 240) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (640, 240) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (640, 240) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (640, 240) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (640, 240) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (640, 240) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (640, 240) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (640, 240) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (640, 240) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (640, 240) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (640, 240) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (640, 240) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (640, 240) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (640, 240) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (640, 240) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (640, 240) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (640, 240) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (640, 240) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (640, 240) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (640, 240) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (640, 240) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (640, 240) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (640, 240) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (640, 240) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (640, 240) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (640, 240) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (640, 240) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (640, 240) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (640, 240) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (640, 240) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (640, 240) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (640, 240) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (640, 240) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (640, 240) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (640, 240) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (640, 240) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (640, 240) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (640, 240) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (640, 240) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (640, 240) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (640, 240) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (640, 240) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (640, 240) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (640, 240) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (640, 240) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (640, 240) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (640, 240) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (640, 240) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (640, 240) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (640, 240) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (640, 240) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (640, 240) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (640, 240) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (640, 240) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (640, 240) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (640, 240) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (640, 240) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (640, 240) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (640, 240) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (640, 240) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (640, 240) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (640, 240) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (640, 240) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (640, 240) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (640, 240) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (640, 240) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (640, 240) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (640, 240) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (640, 240) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (640, 240) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (640, 240) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (640, 240) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (640, 240) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (640, 240) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (640, 240) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (640, 240) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (640, 240) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (640, 240) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (640, 240) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd240;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 45
		if (frame_counter == 7'd45 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (640, 260) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (640, 260) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (640, 260) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (640, 260) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (640, 260) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (640, 260) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (640, 260) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (640, 260) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (640, 260) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (640, 260) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (640, 260) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (640, 260) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (640, 260) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (640, 260) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (640, 260) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (640, 260) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (640, 260) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (640, 260) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (640, 260) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (640, 260) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (640, 260) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (640, 260) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (640, 260) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (640, 260) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (640, 260) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (640, 260) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (640, 260) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (640, 260) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (640, 260) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (640, 260) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (640, 260) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (640, 260) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (640, 260) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (640, 260) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (640, 260) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (640, 260) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (640, 260) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (640, 260) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (640, 260) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (640, 260) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (640, 260) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (640, 260) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (640, 260) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (640, 260) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (640, 260) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (640, 260) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (640, 260) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (640, 260) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (640, 260) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (640, 260) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (640, 260) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (640, 260) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (640, 260) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (640, 260) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (640, 260) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (640, 260) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (640, 260) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (640, 260) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (640, 260) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (640, 260) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (640, 260) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (640, 260) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (640, 260) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (640, 260) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (640, 260) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (640, 260) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (640, 260) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (640, 260) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (640, 260) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (640, 260) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (640, 260) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (640, 260) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (640, 260) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (640, 260) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (640, 260) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (640, 260) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (640, 260) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (640, 260) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (640, 260) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (640, 260) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (640, 260) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (640, 260) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (640, 260) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (640, 260) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (640, 260) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (640, 260) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (640, 260) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (640, 260) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (640, 260) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (640, 260) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (640, 260) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (640, 260) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (640, 260) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (640, 260) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (640, 260) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (640, 260) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (640, 260) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (640, 260) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (640, 260) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (640, 260) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (640, 260) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (640, 260) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (640, 260) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (640, 260) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (640, 260) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (640, 260) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (640, 260) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (640, 260) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (640, 260) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (640, 260) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (640, 260) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (640, 260) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd260;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 46
		if (frame_counter == 7'd46 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (640, 280) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (640, 280) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (640, 280) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (640, 280) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (640, 280) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (640, 280) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (640, 280) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (640, 280) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (640, 280) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (640, 280) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (640, 280) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (640, 280) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (640, 280) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (640, 280) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (640, 280) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (640, 280) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (640, 280) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (640, 280) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (640, 280) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (640, 280) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (640, 280) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (640, 280) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (640, 280) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (640, 280) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (640, 280) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (640, 280) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (640, 280) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (640, 280) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (640, 280) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (640, 280) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (640, 280) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (640, 280) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (640, 280) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (640, 280) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (640, 280) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (640, 280) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (640, 280) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (640, 280) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (640, 280) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (640, 280) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (640, 280) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (640, 280) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (640, 280) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (640, 280) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (640, 280) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (640, 280) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (640, 280) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (640, 280) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (640, 280) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (640, 280) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (640, 280) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (640, 280) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (640, 280) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (640, 280) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (640, 280) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (640, 280) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (640, 280) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (640, 280) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (640, 280) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (640, 280) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (640, 280) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (640, 280) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (640, 280) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (640, 280) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (640, 280) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (640, 280) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (640, 280) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (640, 280) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (640, 280) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (640, 280) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (640, 280) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (640, 280) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (640, 280) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (640, 280) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (640, 280) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (640, 280) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (640, 280) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (640, 280) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (640, 280) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (640, 280) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (640, 280) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (640, 280) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (640, 280) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (640, 280) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (640, 280) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (640, 280) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (640, 280) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (640, 280) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (640, 280) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (640, 280) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (640, 280) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (640, 280) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (640, 280) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (640, 280) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (640, 280) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (640, 280) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (640, 280) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (640, 280) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (640, 280) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (640, 280) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (640, 280) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (640, 280) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (640, 280) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (640, 280) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (640, 280) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (640, 280) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (640, 280) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (640, 280) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (640, 280) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (640, 280) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (640, 280) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (640, 280) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd280;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 47
		if (frame_counter == 7'd47 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (640, 300) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (640, 300) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (640, 300) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (640, 300) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (640, 300) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (640, 300) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (640, 300) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (640, 300) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (640, 300) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (640, 300) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (640, 300) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (640, 300) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (640, 300) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (640, 300) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (640, 300) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (640, 300) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (640, 300) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (640, 300) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (640, 300) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (640, 300) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (640, 300) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (640, 300) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (640, 300) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (640, 300) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (640, 300) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (640, 300) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (640, 300) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (640, 300) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (640, 300) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (640, 300) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (640, 300) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (640, 300) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (640, 300) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (640, 300) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (640, 300) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (640, 300) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (640, 300) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (640, 300) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (640, 300) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (640, 300) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (640, 300) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (640, 300) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (640, 300) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (640, 300) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (640, 300) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (640, 300) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (640, 300) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (640, 300) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (640, 300) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (640, 300) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (640, 300) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (640, 300) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (640, 300) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (640, 300) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (640, 300) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (640, 300) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (640, 300) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (640, 300) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (640, 300) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (640, 300) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (640, 300) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (640, 300) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (640, 300) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (640, 300) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (640, 300) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (640, 300) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (640, 300) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (640, 300) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (640, 300) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (640, 300) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (640, 300) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (640, 300) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (640, 300) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (640, 300) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (640, 300) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (640, 300) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (640, 300) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (640, 300) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (640, 300) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (640, 300) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (640, 300) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (640, 300) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (640, 300) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (640, 300) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (640, 300) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (640, 300) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (640, 300) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (640, 300) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (640, 300) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (640, 300) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (640, 300) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (640, 300) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (640, 300) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (640, 300) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (640, 300) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (640, 300) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (640, 300) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (640, 300) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (640, 300) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (640, 300) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (640, 300) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (640, 300) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (640, 300) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (640, 300) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (640, 300) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (640, 300) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (640, 300) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (640, 300) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (640, 300) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (640, 300) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (640, 300) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (640, 300) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd300;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 48
		if (frame_counter == 7'd48 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (640, 320) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (640, 320) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (640, 320) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (640, 320) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (640, 320) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (640, 320) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (640, 320) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (640, 320) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (640, 320) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (640, 320) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (640, 320) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (640, 320) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (640, 320) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (640, 320) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (640, 320) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (640, 320) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (640, 320) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (640, 320) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (640, 320) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (640, 320) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (640, 320) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (640, 320) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (640, 320) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (640, 320) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (640, 320) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (640, 320) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (640, 320) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (640, 320) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (640, 320) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (640, 320) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (640, 320) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (640, 320) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (640, 320) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (640, 320) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (640, 320) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (640, 320) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (640, 320) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (640, 320) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (640, 320) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (640, 320) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (640, 320) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (640, 320) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (640, 320) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (640, 320) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (640, 320) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (640, 320) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (640, 320) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (640, 320) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (640, 320) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (640, 320) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (640, 320) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (640, 320) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (640, 320) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (640, 320) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (640, 320) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (640, 320) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (640, 320) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (640, 320) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (640, 320) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (640, 320) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (640, 320) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (640, 320) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (640, 320) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (640, 320) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (640, 320) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (640, 320) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (640, 320) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (640, 320) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (640, 320) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (640, 320) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (640, 320) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (640, 320) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (640, 320) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (640, 320) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (640, 320) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (640, 320) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (640, 320) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (640, 320) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (640, 320) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (640, 320) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (640, 320) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (640, 320) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (640, 320) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (640, 320) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (640, 320) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (640, 320) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (640, 320) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (640, 320) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (640, 320) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (640, 320) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (640, 320) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (640, 320) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (640, 320) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (640, 320) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (640, 320) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (640, 320) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (640, 320) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (640, 320) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (640, 320) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (640, 320) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (640, 320) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (640, 320) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (640, 320) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (640, 320) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (640, 320) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (640, 320) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (640, 320) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (640, 320) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (640, 320) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (640, 320) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (640, 320) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (640, 320) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd320;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 49
		if (frame_counter == 7'd49 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (640, 340) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (640, 340) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (640, 340) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (640, 340) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (640, 340) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (640, 340) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (640, 340) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (640, 340) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (640, 340) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (640, 340) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (640, 340) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (640, 340) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (640, 340) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (640, 340) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (640, 340) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (640, 340) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (640, 340) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (640, 340) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (640, 340) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (640, 340) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (640, 340) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (640, 340) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (640, 340) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (640, 340) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (640, 340) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (640, 340) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (640, 340) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (640, 340) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (640, 340) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (640, 340) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (640, 340) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (640, 340) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (640, 340) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (640, 340) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (640, 340) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (640, 340) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (640, 340) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (640, 340) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (640, 340) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (640, 340) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (640, 340) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (640, 340) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (640, 340) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (640, 340) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (640, 340) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (640, 340) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (640, 340) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (640, 340) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (640, 340) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (640, 340) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (640, 340) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (640, 340) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (640, 340) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (640, 340) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (640, 340) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (640, 340) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (640, 340) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (640, 340) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (640, 340) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (640, 340) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (640, 340) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (640, 340) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (640, 340) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (640, 340) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (640, 340) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (640, 340) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (640, 340) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (640, 340) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (640, 340) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (640, 340) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (640, 340) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (640, 340) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (640, 340) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (640, 340) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (640, 340) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (640, 340) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (640, 340) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (640, 340) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (640, 340) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (640, 340) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (640, 340) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (640, 340) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (640, 340) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (640, 340) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (640, 340) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (640, 340) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (640, 340) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (640, 340) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (640, 340) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (640, 340) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (640, 340) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (640, 340) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (640, 340) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (640, 340) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (640, 340) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (640, 340) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (640, 340) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (640, 340) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (640, 340) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (640, 340) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (640, 340) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (640, 340) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (640, 340) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (640, 340) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (640, 340) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (640, 340) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (640, 340) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (640, 340) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (640, 340) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (640, 340) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (640, 340) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (640, 340) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd340;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 50
		if (frame_counter == 7'd50 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (640, 360) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (640, 360) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (640, 360) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (640, 360) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (640, 360) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (640, 360) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (640, 360) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (640, 360) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (640, 360) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (640, 360) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (640, 360) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (640, 360) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (640, 360) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (640, 360) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (640, 360) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (640, 360) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (640, 360) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (640, 360) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (640, 360) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (640, 360) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (640, 360) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (640, 360) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (640, 360) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (640, 360) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (640, 360) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (640, 360) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (640, 360) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (640, 360) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (640, 360) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (640, 360) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (640, 360) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (640, 360) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (640, 360) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (640, 360) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (640, 360) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (640, 360) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (640, 360) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (640, 360) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (640, 360) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (640, 360) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (640, 360) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (640, 360) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (640, 360) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (640, 360) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (640, 360) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (640, 360) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (640, 360) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (640, 360) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (640, 360) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (640, 360) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (640, 360) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (640, 360) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (640, 360) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (640, 360) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (640, 360) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (640, 360) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (640, 360) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (640, 360) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (640, 360) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (640, 360) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (640, 360) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (640, 360) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (640, 360) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (640, 360) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (640, 360) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (640, 360) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (640, 360) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (640, 360) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (640, 360) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (640, 360) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (640, 360) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (640, 360) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (640, 360) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (640, 360) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (640, 360) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (640, 360) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (640, 360) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (640, 360) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (640, 360) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (640, 360) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (640, 360) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (640, 360) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (640, 360) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (640, 360) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (640, 360) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (640, 360) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (640, 360) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (640, 360) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (640, 360) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (640, 360) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (640, 360) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (640, 360) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (640, 360) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (640, 360) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (640, 360) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (640, 360) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (640, 360) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (640, 360) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (640, 360) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (640, 360) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (640, 360) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (640, 360) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (640, 360) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (640, 360) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (640, 360) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (640, 360) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (640, 360) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (640, 360) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (640, 360) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (640, 360) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (640, 360) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (640, 360) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd360;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 51
		if (frame_counter == 7'd51 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (640, 380) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (640, 380) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (640, 380) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (640, 380) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (640, 380) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (640, 380) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (640, 380) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (640, 380) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (640, 380) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (640, 380) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (640, 380) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (640, 380) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (640, 380) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (640, 380) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (640, 380) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (640, 380) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (640, 380) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (640, 380) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (640, 380) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (640, 380) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (640, 380) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (640, 380) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (640, 380) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (640, 380) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (640, 380) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (640, 380) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (640, 380) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (640, 380) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (640, 380) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (640, 380) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (640, 380) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (640, 380) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (640, 380) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (640, 380) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (640, 380) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (640, 380) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (640, 380) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (640, 380) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (640, 380) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (640, 380) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (640, 380) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (640, 380) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (640, 380) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (640, 380) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (640, 380) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (640, 380) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (640, 380) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (640, 380) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (640, 380) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (640, 380) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (640, 380) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (640, 380) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (640, 380) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (640, 380) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (640, 380) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (640, 380) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (640, 380) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (640, 380) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (640, 380) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (640, 380) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (640, 380) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (640, 380) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (640, 380) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (640, 380) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (640, 380) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (640, 380) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (640, 380) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (640, 380) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (640, 380) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (640, 380) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (640, 380) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (640, 380) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (640, 380) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (640, 380) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (640, 380) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (640, 380) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (640, 380) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (640, 380) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (640, 380) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (640, 380) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (640, 380) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (640, 380) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (640, 380) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (640, 380) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (640, 380) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (640, 380) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (640, 380) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (640, 380) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (640, 380) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (640, 380) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (640, 380) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (640, 380) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (640, 380) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (640, 380) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (640, 380) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (640, 380) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (640, 380) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (640, 380) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (640, 380) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (640, 380) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (640, 380) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (640, 380) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (640, 380) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (640, 380) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (640, 380) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (640, 380) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (640, 380) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (640, 380) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (640, 380) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (640, 380) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (640, 380) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (640, 380) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd380;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 52
		if (frame_counter == 7'd52 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (640, 400) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (640, 400) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (640, 400) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (640, 400) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (640, 400) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (640, 400) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (640, 400) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (640, 400) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (640, 400) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (640, 400) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (640, 400) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (640, 400) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (640, 400) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (640, 400) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (640, 400) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (640, 400) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (640, 400) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (640, 400) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (640, 400) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (640, 400) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (640, 400) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (640, 400) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (640, 400) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (640, 400) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (640, 400) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (640, 400) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (640, 400) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (640, 400) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (640, 400) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (640, 400) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (640, 400) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (640, 400) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (640, 400) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (640, 400) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (640, 400) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (640, 400) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (640, 400) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (640, 400) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (640, 400) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (640, 400) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (640, 400) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (640, 400) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (640, 400) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (640, 400) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (640, 400) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (640, 400) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (640, 400) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (640, 400) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (640, 400) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (640, 400) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (640, 400) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (640, 400) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (640, 400) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (640, 400) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (640, 400) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (640, 400) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (640, 400) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (640, 400) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (640, 400) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (640, 400) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (640, 400) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (640, 400) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (640, 400) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (640, 400) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (640, 400) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (640, 400) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (640, 400) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (640, 400) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (640, 400) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (640, 400) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (640, 400) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (640, 400) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (640, 400) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (640, 400) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (640, 400) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (640, 400) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (640, 400) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (640, 400) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (640, 400) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (640, 400) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (640, 400) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (640, 400) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (640, 400) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (640, 400) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (640, 400) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (640, 400) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (640, 400) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (640, 400) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (640, 400) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (640, 400) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (640, 400) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (640, 400) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (640, 400) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (640, 400) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (640, 400) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (640, 400) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (640, 400) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (640, 400) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (640, 400) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (640, 400) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (640, 400) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (640, 400) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (640, 400) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (640, 400) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (640, 400) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (640, 400) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (640, 400) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (640, 400) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (640, 400) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (640, 400) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (640, 400) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (640, 400) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd400;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 53
		if (frame_counter == 7'd53 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (640, 420) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (640, 420) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (640, 420) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (640, 420) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (640, 420) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (640, 420) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (640, 420) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (640, 420) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (640, 420) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (640, 420) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (640, 420) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (640, 420) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (640, 420) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (640, 420) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (640, 420) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (640, 420) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (640, 420) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (640, 420) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (640, 420) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (640, 420) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (640, 420) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (640, 420) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (640, 420) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (640, 420) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (640, 420) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (640, 420) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (640, 420) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (640, 420) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (640, 420) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (640, 420) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (640, 420) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (640, 420) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (640, 420) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (640, 420) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (640, 420) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (640, 420) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (640, 420) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (640, 420) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (640, 420) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (640, 420) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (640, 420) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (640, 420) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (640, 420) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (640, 420) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (640, 420) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (640, 420) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (640, 420) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (640, 420) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (640, 420) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (640, 420) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (640, 420) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (640, 420) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (640, 420) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (640, 420) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (640, 420) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (640, 420) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (640, 420) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (640, 420) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (640, 420) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (640, 420) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (640, 420) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (640, 420) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (640, 420) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (640, 420) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (640, 420) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (640, 420) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (640, 420) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (640, 420) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (640, 420) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (640, 420) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (640, 420) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (640, 420) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (640, 420) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (640, 420) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (640, 420) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (640, 420) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (640, 420) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (640, 420) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (640, 420) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (640, 420) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (640, 420) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (640, 420) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (640, 420) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (640, 420) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (640, 420) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (640, 420) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (640, 420) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (640, 420) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (640, 420) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (640, 420) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (640, 420) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (640, 420) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (640, 420) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (640, 420) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (640, 420) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (640, 420) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (640, 420) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (640, 420) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (640, 420) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (640, 420) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (640, 420) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (640, 420) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (640, 420) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (640, 420) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (640, 420) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (640, 420) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (640, 420) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (640, 420) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (640, 420) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (640, 420) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (640, 420) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (640, 420) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd420;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 54
		if (frame_counter == 7'd54 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (640, 440) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (640, 440) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (640, 440) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (640, 440) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (640, 440) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (640, 440) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (640, 440) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (640, 440) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (640, 440) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (640, 440) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (640, 440) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (640, 440) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (640, 440) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (640, 440) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (640, 440) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (640, 440) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (640, 440) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (640, 440) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (640, 440) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (640, 440) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (640, 440) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (640, 440) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (640, 440) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (640, 440) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (640, 440) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (640, 440) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (640, 440) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (640, 440) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (640, 440) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (640, 440) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (640, 440) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (640, 440) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (640, 440) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (640, 440) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (640, 440) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (640, 440) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (640, 440) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (640, 440) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (640, 440) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (640, 440) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (640, 440) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (640, 440) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (640, 440) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (640, 440) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (640, 440) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (640, 440) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (640, 440) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (640, 440) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (640, 440) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (640, 440) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (640, 440) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (640, 440) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (640, 440) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (640, 440) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (640, 440) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (640, 440) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (640, 440) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (640, 440) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (640, 440) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (640, 440) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (640, 440) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (640, 440) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (640, 440) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (640, 440) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (640, 440) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (640, 440) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (640, 440) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (640, 440) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (640, 440) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (640, 440) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (640, 440) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (640, 440) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (640, 440) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (640, 440) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (640, 440) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (640, 440) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (640, 440) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (640, 440) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (640, 440) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (640, 440) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (640, 440) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (640, 440) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (640, 440) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (640, 440) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (640, 440) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (640, 440) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (640, 440) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (640, 440) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (640, 440) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (640, 440) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (640, 440) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (640, 440) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (640, 440) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (640, 440) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (640, 440) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (640, 440) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (640, 440) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (640, 440) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (640, 440) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (640, 440) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (640, 440) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (640, 440) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (640, 440) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (640, 440) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (640, 440) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (640, 440) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (640, 440) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (640, 440) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (640, 440) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (640, 440) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (640, 440) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (640, 440) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd440;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 55
		if (frame_counter == 7'd55 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (640, 460) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (640, 460) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (640, 460) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (640, 460) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (640, 460) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (640, 460) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (640, 460) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (640, 460) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (640, 460) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (640, 460) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (640, 460) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (640, 460) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (640, 460) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (640, 460) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (640, 460) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (640, 460) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (640, 460) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (640, 460) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (640, 460) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (640, 460) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (640, 460) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (640, 460) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (640, 460) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (640, 460) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (640, 460) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (640, 460) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (640, 460) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (640, 460) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (640, 460) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (640, 460) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (640, 460) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (640, 460) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (640, 460) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (640, 460) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (640, 460) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (640, 460) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (640, 460) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (640, 460) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (640, 460) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (640, 460) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (640, 460) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (640, 460) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (640, 460) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (640, 460) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (640, 460) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (640, 460) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (640, 460) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (640, 460) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (640, 460) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (640, 460) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (640, 460) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (640, 460) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (640, 460) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (640, 460) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (640, 460) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (640, 460) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (640, 460) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (640, 460) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (640, 460) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (640, 460) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (640, 460) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (640, 460) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (640, 460) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (640, 460) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (640, 460) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (640, 460) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (640, 460) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (640, 460) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (640, 460) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (640, 460) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (640, 460) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (640, 460) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (640, 460) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (640, 460) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (640, 460) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (640, 460) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (640, 460) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (640, 460) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (640, 460) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (640, 460) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (640, 460) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (640, 460) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (640, 460) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (640, 460) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (640, 460) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (640, 460) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (640, 460) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (640, 460) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (640, 460) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (640, 460) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (640, 460) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (640, 460) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (640, 460) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (640, 460) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (640, 460) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (640, 460) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (640, 460) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (640, 460) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (640, 460) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (640, 460) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (640, 460) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (640, 460) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (640, 460) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (640, 460) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (640, 460) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (640, 460) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (640, 460) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (640, 460) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (640, 460) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (640, 460) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (640, 460) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (640, 460) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd460;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 56
		if (frame_counter == 7'd56 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (640, 480) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (640, 480) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (640, 480) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (640, 480) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (640, 480) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (640, 480) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (640, 480) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (640, 480) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (640, 480) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (640, 480) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (640, 480) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (640, 480) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (640, 480) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (640, 480) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (640, 480) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (640, 480) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (640, 480) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (640, 480) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (640, 480) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (640, 480) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (640, 480) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (640, 480) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (640, 480) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (640, 480) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (640, 480) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (640, 480) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (640, 480) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (640, 480) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (640, 480) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (640, 480) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (640, 480) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (640, 480) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (640, 480) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (640, 480) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (640, 480) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (640, 480) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (640, 480) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (640, 480) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (640, 480) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (640, 480) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (640, 480) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (640, 480) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (640, 480) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (640, 480) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (640, 480) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (640, 480) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (640, 480) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (640, 480) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (640, 480) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (640, 480) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (640, 480) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (640, 480) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (640, 480) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (640, 480) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (640, 480) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (640, 480) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (640, 480) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (640, 480) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (640, 480) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (640, 480) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (640, 480) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (640, 480) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (640, 480) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (640, 480) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (640, 480) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (640, 480) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (640, 480) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (640, 480) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (640, 480) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (640, 480) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (640, 480) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (640, 480) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (640, 480) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (640, 480) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (640, 480) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (640, 480) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (640, 480) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (640, 480) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (640, 480) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (640, 480) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (640, 480) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (640, 480) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (640, 480) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (640, 480) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (640, 480) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (640, 480) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (640, 480) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (640, 480) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (640, 480) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (640, 480) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (640, 480) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (640, 480) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (640, 480) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (640, 480) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (640, 480) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (640, 480) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (640, 480) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (640, 480) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (640, 480) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (640, 480) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (640, 480) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (640, 480) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (640, 480) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (640, 480) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (640, 480) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (640, 480) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (640, 480) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (640, 480) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (640, 480) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (640, 480) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (640, 480) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (640, 480) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd640;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 57
		if (frame_counter == 7'd57 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (620, 480) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (620, 480) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (620, 480) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (620, 480) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (620, 480) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (620, 480) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (620, 480) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (620, 480) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (620, 480) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (620, 480) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (620, 480) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (620, 480) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (620, 480) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (620, 480) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (620, 480) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (620, 480) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (620, 480) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (620, 480) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (620, 480) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (620, 480) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (620, 480) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (620, 480) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (620, 480) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (620, 480) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (620, 480) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (620, 480) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (620, 480) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (620, 480) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (620, 480) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (620, 480) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (620, 480) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (620, 480) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (620, 480) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (620, 480) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (620, 480) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (620, 480) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (620, 480) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (620, 480) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (620, 480) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (620, 480) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (620, 480) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (620, 480) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (620, 480) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (620, 480) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (620, 480) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (620, 480) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (620, 480) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (620, 480) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (620, 480) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (620, 480) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (620, 480) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (620, 480) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (620, 480) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (620, 480) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (620, 480) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (620, 480) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (620, 480) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (620, 480) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (620, 480) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (620, 480) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (620, 480) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (620, 480) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (620, 480) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (620, 480) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (620, 480) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (620, 480) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (620, 480) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (620, 480) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (620, 480) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (620, 480) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (620, 480) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (620, 480) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (620, 480) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (620, 480) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (620, 480) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (620, 480) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (620, 480) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (620, 480) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (620, 480) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (620, 480) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (620, 480) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (620, 480) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (620, 480) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (620, 480) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (620, 480) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (620, 480) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (620, 480) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (620, 480) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (620, 480) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (620, 480) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (620, 480) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (620, 480) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (620, 480) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (620, 480) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (620, 480) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (620, 480) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (620, 480) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (620, 480) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (620, 480) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (620, 480) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (620, 480) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (620, 480) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (620, 480) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (620, 480) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (620, 480) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (620, 480) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (620, 480) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (620, 480) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (620, 480) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (620, 480) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (620, 480) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (620, 480) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd620;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 58
		if (frame_counter == 7'd58 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (600, 480) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (600, 480) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (600, 480) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (600, 480) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (600, 480) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (600, 480) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (600, 480) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (600, 480) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (600, 480) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (600, 480) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (600, 480) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (600, 480) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (600, 480) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (600, 480) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (600, 480) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (600, 480) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (600, 480) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (600, 480) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (600, 480) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (600, 480) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (600, 480) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (600, 480) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (600, 480) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (600, 480) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (600, 480) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (600, 480) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (600, 480) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (600, 480) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (600, 480) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (600, 480) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (600, 480) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (600, 480) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (600, 480) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (600, 480) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (600, 480) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (600, 480) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (600, 480) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (600, 480) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (600, 480) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (600, 480) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (600, 480) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (600, 480) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (600, 480) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (600, 480) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (600, 480) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (600, 480) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (600, 480) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (600, 480) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (600, 480) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (600, 480) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (600, 480) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (600, 480) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (600, 480) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (600, 480) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (600, 480) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (600, 480) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (600, 480) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (600, 480) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (600, 480) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (600, 480) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (600, 480) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (600, 480) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (600, 480) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (600, 480) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (600, 480) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (600, 480) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (600, 480) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (600, 480) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (600, 480) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (600, 480) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (600, 480) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (600, 480) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (600, 480) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (600, 480) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (600, 480) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (600, 480) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (600, 480) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (600, 480) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (600, 480) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (600, 480) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (600, 480) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (600, 480) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (600, 480) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (600, 480) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (600, 480) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (600, 480) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (600, 480) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (600, 480) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (600, 480) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (600, 480) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (600, 480) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (600, 480) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (600, 480) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (600, 480) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (600, 480) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (600, 480) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (600, 480) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (600, 480) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (600, 480) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (600, 480) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (600, 480) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (600, 480) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (600, 480) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (600, 480) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (600, 480) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (600, 480) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (600, 480) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (600, 480) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (600, 480) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (600, 480) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (600, 480) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (600, 480) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd600;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 59
		if (frame_counter == 7'd59 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (580, 480) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (580, 480) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (580, 480) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (580, 480) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (580, 480) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (580, 480) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (580, 480) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (580, 480) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (580, 480) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (580, 480) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (580, 480) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (580, 480) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (580, 480) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (580, 480) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (580, 480) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (580, 480) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (580, 480) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (580, 480) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (580, 480) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (580, 480) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (580, 480) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (580, 480) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (580, 480) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (580, 480) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (580, 480) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (580, 480) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (580, 480) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (580, 480) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (580, 480) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (580, 480) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (580, 480) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (580, 480) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (580, 480) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (580, 480) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (580, 480) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (580, 480) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (580, 480) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (580, 480) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (580, 480) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (580, 480) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (580, 480) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (580, 480) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (580, 480) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (580, 480) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (580, 480) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (580, 480) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (580, 480) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (580, 480) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (580, 480) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (580, 480) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (580, 480) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (580, 480) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (580, 480) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (580, 480) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (580, 480) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (580, 480) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (580, 480) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (580, 480) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (580, 480) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (580, 480) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (580, 480) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (580, 480) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (580, 480) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (580, 480) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (580, 480) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (580, 480) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (580, 480) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (580, 480) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (580, 480) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (580, 480) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (580, 480) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (580, 480) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (580, 480) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (580, 480) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (580, 480) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (580, 480) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (580, 480) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (580, 480) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (580, 480) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (580, 480) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (580, 480) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (580, 480) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (580, 480) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (580, 480) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (580, 480) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (580, 480) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (580, 480) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (580, 480) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (580, 480) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (580, 480) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (580, 480) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (580, 480) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (580, 480) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (580, 480) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (580, 480) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (580, 480) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (580, 480) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (580, 480) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (580, 480) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (580, 480) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (580, 480) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (580, 480) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (580, 480) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (580, 480) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (580, 480) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (580, 480) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (580, 480) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (580, 480) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (580, 480) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (580, 480) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (580, 480) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (580, 480) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd580;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 60
		if (frame_counter == 7'd60 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (560, 480) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (560, 480) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (560, 480) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (560, 480) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (560, 480) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (560, 480) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (560, 480) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (560, 480) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (560, 480) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (560, 480) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (560, 480) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (560, 480) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (560, 480) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (560, 480) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (560, 480) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (560, 480) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (560, 480) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (560, 480) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (560, 480) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (560, 480) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (560, 480) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (560, 480) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (560, 480) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (560, 480) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (560, 480) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (560, 480) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (560, 480) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (560, 480) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (560, 480) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (560, 480) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (560, 480) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (560, 480) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (560, 480) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (560, 480) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (560, 480) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (560, 480) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (560, 480) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (560, 480) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (560, 480) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (560, 480) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (560, 480) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (560, 480) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (560, 480) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (560, 480) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (560, 480) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (560, 480) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (560, 480) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (560, 480) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (560, 480) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (560, 480) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (560, 480) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (560, 480) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (560, 480) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (560, 480) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (560, 480) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (560, 480) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (560, 480) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (560, 480) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (560, 480) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (560, 480) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (560, 480) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (560, 480) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (560, 480) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (560, 480) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (560, 480) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (560, 480) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (560, 480) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (560, 480) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (560, 480) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (560, 480) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (560, 480) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (560, 480) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (560, 480) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (560, 480) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (560, 480) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (560, 480) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (560, 480) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (560, 480) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (560, 480) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (560, 480) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (560, 480) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (560, 480) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (560, 480) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (560, 480) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (560, 480) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (560, 480) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (560, 480) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (560, 480) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (560, 480) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (560, 480) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (560, 480) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (560, 480) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (560, 480) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (560, 480) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (560, 480) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (560, 480) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (560, 480) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (560, 480) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (560, 480) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (560, 480) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (560, 480) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (560, 480) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (560, 480) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (560, 480) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (560, 480) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (560, 480) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (560, 480) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (560, 480) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (560, 480) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (560, 480) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (560, 480) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (560, 480) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd560;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 61
		if (frame_counter == 7'd61 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (540, 480) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (540, 480) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (540, 480) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (540, 480) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (540, 480) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (540, 480) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (540, 480) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (540, 480) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (540, 480) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (540, 480) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (540, 480) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (540, 480) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (540, 480) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (540, 480) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (540, 480) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (540, 480) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (540, 480) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (540, 480) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (540, 480) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (540, 480) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (540, 480) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (540, 480) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (540, 480) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (540, 480) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (540, 480) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (540, 480) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (540, 480) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (540, 480) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (540, 480) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (540, 480) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (540, 480) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (540, 480) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (540, 480) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (540, 480) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (540, 480) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (540, 480) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (540, 480) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (540, 480) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (540, 480) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (540, 480) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (540, 480) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (540, 480) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (540, 480) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (540, 480) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (540, 480) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (540, 480) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (540, 480) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (540, 480) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (540, 480) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (540, 480) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (540, 480) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (540, 480) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (540, 480) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (540, 480) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (540, 480) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (540, 480) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (540, 480) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (540, 480) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (540, 480) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (540, 480) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (540, 480) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (540, 480) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (540, 480) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (540, 480) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (540, 480) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (540, 480) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (540, 480) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (540, 480) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (540, 480) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (540, 480) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (540, 480) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (540, 480) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (540, 480) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (540, 480) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (540, 480) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (540, 480) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (540, 480) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (540, 480) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (540, 480) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (540, 480) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (540, 480) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (540, 480) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (540, 480) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (540, 480) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (540, 480) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (540, 480) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (540, 480) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (540, 480) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (540, 480) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (540, 480) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (540, 480) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (540, 480) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (540, 480) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (540, 480) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (540, 480) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (540, 480) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (540, 480) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (540, 480) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (540, 480) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (540, 480) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (540, 480) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (540, 480) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (540, 480) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (540, 480) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (540, 480) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (540, 480) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (540, 480) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (540, 480) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (540, 480) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (540, 480) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (540, 480) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (540, 480) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd540;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 62
		if (frame_counter == 7'd62 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (520, 480) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (520, 480) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (520, 480) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (520, 480) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (520, 480) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (520, 480) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (520, 480) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (520, 480) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (520, 480) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (520, 480) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (520, 480) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (520, 480) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (520, 480) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (520, 480) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (520, 480) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (520, 480) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (520, 480) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (520, 480) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (520, 480) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (520, 480) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (520, 480) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (520, 480) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (520, 480) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (520, 480) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (520, 480) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (520, 480) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (520, 480) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (520, 480) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (520, 480) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (520, 480) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (520, 480) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (520, 480) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (520, 480) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (520, 480) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (520, 480) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (520, 480) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (520, 480) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (520, 480) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (520, 480) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (520, 480) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (520, 480) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (520, 480) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (520, 480) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (520, 480) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (520, 480) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (520, 480) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (520, 480) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (520, 480) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (520, 480) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (520, 480) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (520, 480) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (520, 480) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (520, 480) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (520, 480) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (520, 480) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (520, 480) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (520, 480) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (520, 480) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (520, 480) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (520, 480) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (520, 480) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (520, 480) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (520, 480) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (520, 480) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (520, 480) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (520, 480) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (520, 480) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (520, 480) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (520, 480) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (520, 480) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (520, 480) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (520, 480) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (520, 480) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (520, 480) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (520, 480) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (520, 480) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (520, 480) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (520, 480) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (520, 480) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (520, 480) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (520, 480) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (520, 480) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (520, 480) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (520, 480) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (520, 480) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (520, 480) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (520, 480) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (520, 480) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (520, 480) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (520, 480) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (520, 480) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (520, 480) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (520, 480) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (520, 480) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (520, 480) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (520, 480) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (520, 480) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (520, 480) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (520, 480) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (520, 480) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (520, 480) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (520, 480) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (520, 480) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (520, 480) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (520, 480) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (520, 480) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (520, 480) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (520, 480) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (520, 480) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (520, 480) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (520, 480) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (520, 480) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd520;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 63
		if (frame_counter == 7'd63 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (500, 480) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (500, 480) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (500, 480) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (500, 480) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (500, 480) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (500, 480) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (500, 480) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (500, 480) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (500, 480) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (500, 480) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (500, 480) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (500, 480) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (500, 480) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (500, 480) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (500, 480) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (500, 480) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (500, 480) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (500, 480) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (500, 480) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (500, 480) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (500, 480) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (500, 480) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (500, 480) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (500, 480) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (500, 480) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (500, 480) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (500, 480) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (500, 480) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (500, 480) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (500, 480) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (500, 480) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (500, 480) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (500, 480) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (500, 480) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (500, 480) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (500, 480) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (500, 480) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (500, 480) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (500, 480) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (500, 480) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (500, 480) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (500, 480) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (500, 480) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (500, 480) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (500, 480) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (500, 480) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (500, 480) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (500, 480) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (500, 480) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (500, 480) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (500, 480) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (500, 480) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (500, 480) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (500, 480) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (500, 480) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (500, 480) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (500, 480) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (500, 480) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (500, 480) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (500, 480) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (500, 480) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (500, 480) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (500, 480) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (500, 480) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (500, 480) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (500, 480) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (500, 480) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (500, 480) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (500, 480) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (500, 480) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (500, 480) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (500, 480) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (500, 480) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (500, 480) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (500, 480) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (500, 480) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (500, 480) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (500, 480) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (500, 480) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (500, 480) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (500, 480) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (500, 480) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (500, 480) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (500, 480) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (500, 480) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (500, 480) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (500, 480) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (500, 480) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (500, 480) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (500, 480) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (500, 480) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (500, 480) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (500, 480) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (500, 480) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (500, 480) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (500, 480) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (500, 480) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (500, 480) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (500, 480) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (500, 480) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (500, 480) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (500, 480) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (500, 480) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (500, 480) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (500, 480) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (500, 480) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (500, 480) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (500, 480) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (500, 480) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (500, 480) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (500, 480) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (500, 480) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd500;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 64
		if (frame_counter == 7'd64 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (480, 480) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (480, 480) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (480, 480) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (480, 480) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (480, 480) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (480, 480) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (480, 480) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (480, 480) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (480, 480) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (480, 480) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (480, 480) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (480, 480) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (480, 480) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (480, 480) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (480, 480) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (480, 480) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (480, 480) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (480, 480) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (480, 480) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (480, 480) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (480, 480) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (480, 480) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (480, 480) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (480, 480) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (480, 480) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (480, 480) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (480, 480) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (480, 480) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (480, 480) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (480, 480) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (480, 480) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (480, 480) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (480, 480) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (480, 480) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (480, 480) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (480, 480) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (480, 480) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (480, 480) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (480, 480) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (480, 480) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (480, 480) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (480, 480) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (480, 480) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (480, 480) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (480, 480) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (480, 480) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (480, 480) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (480, 480) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (480, 480) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (480, 480) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (480, 480) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (480, 480) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (480, 480) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (480, 480) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (480, 480) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (480, 480) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (480, 480) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (480, 480) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (480, 480) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (480, 480) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (480, 480) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (480, 480) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (480, 480) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (480, 480) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (480, 480) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (480, 480) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (480, 480) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (480, 480) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (480, 480) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (480, 480) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (480, 480) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (480, 480) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (480, 480) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (480, 480) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (480, 480) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (480, 480) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (480, 480) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (480, 480) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (480, 480) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (480, 480) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (480, 480) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (480, 480) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (480, 480) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (480, 480) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (480, 480) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (480, 480) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (480, 480) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (480, 480) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (480, 480) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (480, 480) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (480, 480) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (480, 480) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (480, 480) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (480, 480) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (480, 480) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (480, 480) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (480, 480) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (480, 480) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (480, 480) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (480, 480) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (480, 480) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (480, 480) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (480, 480) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (480, 480) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (480, 480) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (480, 480) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (480, 480) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (480, 480) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (480, 480) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (480, 480) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (480, 480) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (480, 480) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd480;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 65
		if (frame_counter == 7'd65 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (460, 480) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (460, 480) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (460, 480) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (460, 480) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (460, 480) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (460, 480) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (460, 480) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (460, 480) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (460, 480) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (460, 480) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (460, 480) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (460, 480) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (460, 480) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (460, 480) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (460, 480) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (460, 480) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (460, 480) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (460, 480) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (460, 480) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (460, 480) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (460, 480) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (460, 480) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (460, 480) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (460, 480) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (460, 480) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (460, 480) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (460, 480) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (460, 480) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (460, 480) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (460, 480) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (460, 480) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (460, 480) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (460, 480) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (460, 480) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (460, 480) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (460, 480) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (460, 480) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (460, 480) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (460, 480) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (460, 480) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (460, 480) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (460, 480) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (460, 480) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (460, 480) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (460, 480) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (460, 480) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (460, 480) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (460, 480) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (460, 480) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (460, 480) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (460, 480) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (460, 480) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (460, 480) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (460, 480) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (460, 480) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (460, 480) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (460, 480) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (460, 480) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (460, 480) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (460, 480) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (460, 480) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (460, 480) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (460, 480) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (460, 480) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (460, 480) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (460, 480) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (460, 480) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (460, 480) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (460, 480) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (460, 480) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (460, 480) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (460, 480) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (460, 480) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (460, 480) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (460, 480) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (460, 480) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (460, 480) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (460, 480) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (460, 480) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (460, 480) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (460, 480) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (460, 480) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (460, 480) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (460, 480) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (460, 480) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (460, 480) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (460, 480) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (460, 480) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (460, 480) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (460, 480) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (460, 480) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (460, 480) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (460, 480) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (460, 480) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (460, 480) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (460, 480) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (460, 480) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (460, 480) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (460, 480) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (460, 480) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (460, 480) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (460, 480) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (460, 480) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (460, 480) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (460, 480) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (460, 480) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (460, 480) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (460, 480) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (460, 480) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (460, 480) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (460, 480) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (460, 480) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd460;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 66
		if (frame_counter == 7'd66 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (440, 480) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (440, 480) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (440, 480) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (440, 480) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (440, 480) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (440, 480) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (440, 480) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (440, 480) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (440, 480) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (440, 480) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (440, 480) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (440, 480) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (440, 480) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (440, 480) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (440, 480) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (440, 480) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (440, 480) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (440, 480) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (440, 480) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (440, 480) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (440, 480) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (440, 480) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (440, 480) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (440, 480) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (440, 480) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (440, 480) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (440, 480) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (440, 480) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (440, 480) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (440, 480) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (440, 480) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (440, 480) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (440, 480) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (440, 480) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (440, 480) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (440, 480) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (440, 480) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (440, 480) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (440, 480) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (440, 480) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (440, 480) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (440, 480) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (440, 480) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (440, 480) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (440, 480) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (440, 480) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (440, 480) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (440, 480) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (440, 480) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (440, 480) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (440, 480) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (440, 480) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (440, 480) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (440, 480) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (440, 480) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (440, 480) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (440, 480) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (440, 480) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (440, 480) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (440, 480) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (440, 480) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (440, 480) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (440, 480) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (440, 480) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (440, 480) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (440, 480) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (440, 480) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (440, 480) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (440, 480) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (440, 480) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (440, 480) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (440, 480) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (440, 480) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (440, 480) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (440, 480) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (440, 480) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (440, 480) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (440, 480) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (440, 480) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (440, 480) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (440, 480) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (440, 480) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (440, 480) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (440, 480) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (440, 480) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (440, 480) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (440, 480) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (440, 480) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (440, 480) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (440, 480) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (440, 480) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (440, 480) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (440, 480) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (440, 480) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (440, 480) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (440, 480) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (440, 480) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (440, 480) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (440, 480) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (440, 480) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (440, 480) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (440, 480) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (440, 480) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (440, 480) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (440, 480) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (440, 480) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (440, 480) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (440, 480) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (440, 480) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (440, 480) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (440, 480) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (440, 480) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd440;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 67
		if (frame_counter == 7'd67 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (420, 480) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (420, 480) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (420, 480) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (420, 480) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (420, 480) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (420, 480) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (420, 480) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (420, 480) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (420, 480) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (420, 480) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (420, 480) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (420, 480) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (420, 480) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (420, 480) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (420, 480) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (420, 480) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (420, 480) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (420, 480) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (420, 480) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (420, 480) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (420, 480) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (420, 480) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (420, 480) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (420, 480) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (420, 480) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (420, 480) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (420, 480) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (420, 480) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (420, 480) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (420, 480) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (420, 480) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (420, 480) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (420, 480) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (420, 480) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (420, 480) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (420, 480) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (420, 480) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (420, 480) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (420, 480) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (420, 480) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (420, 480) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (420, 480) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (420, 480) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (420, 480) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (420, 480) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (420, 480) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (420, 480) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (420, 480) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (420, 480) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (420, 480) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (420, 480) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (420, 480) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (420, 480) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (420, 480) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (420, 480) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (420, 480) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (420, 480) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (420, 480) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (420, 480) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (420, 480) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (420, 480) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (420, 480) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (420, 480) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (420, 480) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (420, 480) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (420, 480) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (420, 480) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (420, 480) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (420, 480) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (420, 480) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (420, 480) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (420, 480) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (420, 480) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (420, 480) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (420, 480) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (420, 480) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (420, 480) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (420, 480) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (420, 480) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (420, 480) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (420, 480) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (420, 480) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (420, 480) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (420, 480) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (420, 480) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (420, 480) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (420, 480) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (420, 480) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (420, 480) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (420, 480) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (420, 480) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (420, 480) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (420, 480) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (420, 480) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (420, 480) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (420, 480) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (420, 480) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (420, 480) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (420, 480) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (420, 480) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (420, 480) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (420, 480) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (420, 480) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (420, 480) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (420, 480) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (420, 480) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (420, 480) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (420, 480) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (420, 480) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (420, 480) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (420, 480) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (420, 480) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd420;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 68
		if (frame_counter == 7'd68 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (400, 480) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (400, 480) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (400, 480) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (400, 480) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (400, 480) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (400, 480) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (400, 480) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (400, 480) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (400, 480) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (400, 480) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (400, 480) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (400, 480) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (400, 480) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (400, 480) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (400, 480) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (400, 480) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (400, 480) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (400, 480) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (400, 480) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (400, 480) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (400, 480) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (400, 480) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (400, 480) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (400, 480) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (400, 480) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (400, 480) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (400, 480) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (400, 480) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (400, 480) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (400, 480) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (400, 480) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (400, 480) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (400, 480) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (400, 480) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (400, 480) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (400, 480) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (400, 480) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (400, 480) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (400, 480) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (400, 480) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (400, 480) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (400, 480) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (400, 480) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (400, 480) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (400, 480) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (400, 480) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (400, 480) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (400, 480) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (400, 480) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (400, 480) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (400, 480) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (400, 480) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (400, 480) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (400, 480) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (400, 480) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (400, 480) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (400, 480) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (400, 480) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (400, 480) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (400, 480) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (400, 480) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (400, 480) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (400, 480) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (400, 480) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (400, 480) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (400, 480) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (400, 480) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (400, 480) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (400, 480) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (400, 480) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (400, 480) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (400, 480) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (400, 480) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (400, 480) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (400, 480) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (400, 480) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (400, 480) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (400, 480) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (400, 480) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (400, 480) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (400, 480) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (400, 480) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (400, 480) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (400, 480) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (400, 480) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (400, 480) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (400, 480) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (400, 480) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (400, 480) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (400, 480) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (400, 480) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (400, 480) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (400, 480) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (400, 480) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (400, 480) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (400, 480) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (400, 480) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (400, 480) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (400, 480) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (400, 480) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (400, 480) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (400, 480) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (400, 480) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (400, 480) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (400, 480) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (400, 480) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (400, 480) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (400, 480) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (400, 480) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (400, 480) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (400, 480) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (400, 480) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd400;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 69
		if (frame_counter == 7'd69 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (380, 480) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (380, 480) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (380, 480) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (380, 480) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (380, 480) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (380, 480) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (380, 480) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (380, 480) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (380, 480) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (380, 480) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (380, 480) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (380, 480) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (380, 480) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (380, 480) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (380, 480) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (380, 480) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (380, 480) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (380, 480) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (380, 480) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (380, 480) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (380, 480) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (380, 480) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (380, 480) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (380, 480) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (380, 480) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (380, 480) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (380, 480) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (380, 480) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (380, 480) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (380, 480) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (380, 480) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (380, 480) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (380, 480) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (380, 480) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (380, 480) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (380, 480) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (380, 480) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (380, 480) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (380, 480) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (380, 480) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (380, 480) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (380, 480) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (380, 480) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (380, 480) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (380, 480) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (380, 480) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (380, 480) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (380, 480) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (380, 480) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (380, 480) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (380, 480) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (380, 480) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (380, 480) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (380, 480) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (380, 480) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (380, 480) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (380, 480) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (380, 480) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (380, 480) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (380, 480) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (380, 480) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (380, 480) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (380, 480) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (380, 480) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (380, 480) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (380, 480) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (380, 480) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (380, 480) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (380, 480) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (380, 480) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (380, 480) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (380, 480) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (380, 480) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (380, 480) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (380, 480) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (380, 480) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (380, 480) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (380, 480) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (380, 480) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (380, 480) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (380, 480) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (380, 480) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (380, 480) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (380, 480) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (380, 480) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (380, 480) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (380, 480) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (380, 480) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (380, 480) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (380, 480) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (380, 480) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (380, 480) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (380, 480) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (380, 480) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (380, 480) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (380, 480) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (380, 480) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (380, 480) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (380, 480) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (380, 480) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (380, 480) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (380, 480) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (380, 480) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (380, 480) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (380, 480) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (380, 480) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (380, 480) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (380, 480) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (380, 480) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (380, 480) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (380, 480) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (380, 480) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd380;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 70
		if (frame_counter == 7'd70 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (360, 480) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (360, 480) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (360, 480) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (360, 480) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (360, 480) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (360, 480) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (360, 480) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (360, 480) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (360, 480) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (360, 480) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (360, 480) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (360, 480) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (360, 480) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (360, 480) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (360, 480) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (360, 480) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (360, 480) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (360, 480) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (360, 480) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (360, 480) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (360, 480) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (360, 480) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (360, 480) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (360, 480) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (360, 480) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (360, 480) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (360, 480) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (360, 480) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (360, 480) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (360, 480) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (360, 480) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (360, 480) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (360, 480) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (360, 480) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (360, 480) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (360, 480) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (360, 480) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (360, 480) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (360, 480) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (360, 480) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (360, 480) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (360, 480) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (360, 480) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (360, 480) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (360, 480) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (360, 480) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (360, 480) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (360, 480) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (360, 480) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (360, 480) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (360, 480) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (360, 480) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (360, 480) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (360, 480) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (360, 480) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (360, 480) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (360, 480) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (360, 480) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (360, 480) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (360, 480) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (360, 480) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (360, 480) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (360, 480) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (360, 480) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (360, 480) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (360, 480) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (360, 480) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (360, 480) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (360, 480) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (360, 480) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (360, 480) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (360, 480) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (360, 480) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (360, 480) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (360, 480) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (360, 480) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (360, 480) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (360, 480) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (360, 480) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (360, 480) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (360, 480) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (360, 480) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (360, 480) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (360, 480) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (360, 480) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (360, 480) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (360, 480) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (360, 480) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (360, 480) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (360, 480) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (360, 480) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (360, 480) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (360, 480) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (360, 480) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (360, 480) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (360, 480) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (360, 480) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (360, 480) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (360, 480) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (360, 480) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (360, 480) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (360, 480) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (360, 480) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (360, 480) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (360, 480) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (360, 480) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (360, 480) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (360, 480) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (360, 480) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (360, 480) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (360, 480) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (360, 480) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd360;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 71
		if (frame_counter == 7'd71 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (340, 480) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (340, 480) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (340, 480) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (340, 480) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (340, 480) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (340, 480) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (340, 480) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (340, 480) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (340, 480) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (340, 480) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (340, 480) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (340, 480) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (340, 480) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (340, 480) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (340, 480) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (340, 480) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (340, 480) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (340, 480) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (340, 480) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (340, 480) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (340, 480) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (340, 480) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (340, 480) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (340, 480) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (340, 480) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (340, 480) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (340, 480) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (340, 480) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (340, 480) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (340, 480) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (340, 480) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (340, 480) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (340, 480) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (340, 480) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (340, 480) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (340, 480) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (340, 480) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (340, 480) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (340, 480) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (340, 480) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (340, 480) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (340, 480) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (340, 480) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (340, 480) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (340, 480) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (340, 480) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (340, 480) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (340, 480) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (340, 480) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (340, 480) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (340, 480) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (340, 480) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (340, 480) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (340, 480) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (340, 480) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (340, 480) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (340, 480) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (340, 480) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (340, 480) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (340, 480) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (340, 480) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (340, 480) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (340, 480) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (340, 480) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (340, 480) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (340, 480) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (340, 480) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (340, 480) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (340, 480) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (340, 480) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (340, 480) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (340, 480) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (340, 480) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (340, 480) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (340, 480) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (340, 480) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (340, 480) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (340, 480) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (340, 480) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (340, 480) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (340, 480) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (340, 480) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (340, 480) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (340, 480) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (340, 480) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (340, 480) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (340, 480) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (340, 480) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (340, 480) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (340, 480) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (340, 480) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (340, 480) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (340, 480) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (340, 480) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (340, 480) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (340, 480) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (340, 480) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (340, 480) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (340, 480) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (340, 480) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (340, 480) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (340, 480) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (340, 480) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (340, 480) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (340, 480) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (340, 480) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (340, 480) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (340, 480) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (340, 480) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (340, 480) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (340, 480) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (340, 480) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd340;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 72
		if (frame_counter == 7'd72 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (320, 480) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (320, 480) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (320, 480) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (320, 480) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (320, 480) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (320, 480) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (320, 480) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (320, 480) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (320, 480) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (320, 480) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (320, 480) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (320, 480) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (320, 480) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (320, 480) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (320, 480) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (320, 480) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (320, 480) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (320, 480) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (320, 480) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (320, 480) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (320, 480) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (320, 480) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (320, 480) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (320, 480) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (320, 480) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (320, 480) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (320, 480) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (320, 480) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (320, 480) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (320, 480) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (320, 480) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (320, 480) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (320, 480) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (320, 480) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (320, 480) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (320, 480) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (320, 480) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (320, 480) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (320, 480) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (320, 480) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (320, 480) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (320, 480) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (320, 480) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (320, 480) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (320, 480) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (320, 480) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (320, 480) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (320, 480) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (320, 480) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (320, 480) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (320, 480) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (320, 480) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (320, 480) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (320, 480) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (320, 480) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (320, 480) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (320, 480) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (320, 480) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (320, 480) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (320, 480) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (320, 480) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (320, 480) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (320, 480) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (320, 480) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (320, 480) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (320, 480) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (320, 480) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (320, 480) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (320, 480) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (320, 480) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (320, 480) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (320, 480) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (320, 480) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (320, 480) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (320, 480) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (320, 480) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (320, 480) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (320, 480) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (320, 480) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (320, 480) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (320, 480) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (320, 480) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (320, 480) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (320, 480) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (320, 480) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (320, 480) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (320, 480) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (320, 480) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (320, 480) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (320, 480) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (320, 480) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (320, 480) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (320, 480) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (320, 480) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (320, 480) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (320, 480) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (320, 480) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (320, 480) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (320, 480) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (320, 480) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (320, 480) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (320, 480) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (320, 480) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (320, 480) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (320, 480) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (320, 480) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (320, 480) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (320, 480) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (320, 480) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (320, 480) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (320, 480) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (320, 480) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd320;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 73
		if (frame_counter == 7'd73 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (300, 480) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (300, 480) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (300, 480) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (300, 480) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (300, 480) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (300, 480) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (300, 480) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (300, 480) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (300, 480) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (300, 480) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (300, 480) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (300, 480) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (300, 480) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (300, 480) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (300, 480) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (300, 480) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (300, 480) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (300, 480) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (300, 480) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (300, 480) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (300, 480) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (300, 480) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (300, 480) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (300, 480) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (300, 480) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (300, 480) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (300, 480) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (300, 480) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (300, 480) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (300, 480) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (300, 480) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (300, 480) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (300, 480) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (300, 480) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (300, 480) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (300, 480) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (300, 480) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (300, 480) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (300, 480) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (300, 480) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (300, 480) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (300, 480) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (300, 480) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (300, 480) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (300, 480) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (300, 480) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (300, 480) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (300, 480) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (300, 480) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (300, 480) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (300, 480) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (300, 480) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (300, 480) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (300, 480) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (300, 480) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (300, 480) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (300, 480) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (300, 480) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (300, 480) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (300, 480) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (300, 480) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (300, 480) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (300, 480) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (300, 480) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (300, 480) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (300, 480) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (300, 480) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (300, 480) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (300, 480) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (300, 480) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (300, 480) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (300, 480) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (300, 480) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (300, 480) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (300, 480) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (300, 480) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (300, 480) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (300, 480) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (300, 480) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (300, 480) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (300, 480) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (300, 480) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (300, 480) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (300, 480) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (300, 480) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (300, 480) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (300, 480) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (300, 480) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (300, 480) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (300, 480) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (300, 480) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (300, 480) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (300, 480) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (300, 480) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (300, 480) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (300, 480) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (300, 480) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (300, 480) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (300, 480) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (300, 480) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (300, 480) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (300, 480) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (300, 480) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (300, 480) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (300, 480) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (300, 480) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (300, 480) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (300, 480) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (300, 480) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (300, 480) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (300, 480) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (300, 480) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd300;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 74
		if (frame_counter == 7'd74 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (280, 480) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (280, 480) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (280, 480) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (280, 480) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (280, 480) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (280, 480) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (280, 480) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (280, 480) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (280, 480) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (280, 480) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (280, 480) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (280, 480) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (280, 480) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (280, 480) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (280, 480) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (280, 480) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (280, 480) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (280, 480) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (280, 480) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (280, 480) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (280, 480) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (280, 480) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (280, 480) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (280, 480) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (280, 480) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (280, 480) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (280, 480) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (280, 480) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (280, 480) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (280, 480) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (280, 480) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (280, 480) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (280, 480) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (280, 480) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (280, 480) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (280, 480) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (280, 480) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (280, 480) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (280, 480) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (280, 480) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (280, 480) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (280, 480) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (280, 480) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (280, 480) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (280, 480) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (280, 480) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (280, 480) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (280, 480) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (280, 480) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (280, 480) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (280, 480) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (280, 480) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (280, 480) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (280, 480) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (280, 480) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (280, 480) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (280, 480) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (280, 480) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (280, 480) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (280, 480) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (280, 480) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (280, 480) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (280, 480) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (280, 480) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (280, 480) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (280, 480) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (280, 480) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (280, 480) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (280, 480) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (280, 480) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (280, 480) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (280, 480) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (280, 480) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (280, 480) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (280, 480) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (280, 480) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (280, 480) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (280, 480) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (280, 480) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (280, 480) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (280, 480) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (280, 480) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (280, 480) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (280, 480) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (280, 480) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (280, 480) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (280, 480) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (280, 480) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (280, 480) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (280, 480) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (280, 480) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (280, 480) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (280, 480) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (280, 480) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (280, 480) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (280, 480) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (280, 480) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (280, 480) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (280, 480) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (280, 480) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (280, 480) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (280, 480) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (280, 480) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (280, 480) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (280, 480) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (280, 480) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (280, 480) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (280, 480) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (280, 480) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (280, 480) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (280, 480) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (280, 480) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd280;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 75
		if (frame_counter == 7'd75 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (260, 480) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (260, 480) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (260, 480) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (260, 480) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (260, 480) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (260, 480) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (260, 480) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (260, 480) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (260, 480) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (260, 480) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (260, 480) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (260, 480) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (260, 480) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (260, 480) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (260, 480) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (260, 480) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (260, 480) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (260, 480) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (260, 480) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (260, 480) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (260, 480) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (260, 480) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (260, 480) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (260, 480) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (260, 480) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (260, 480) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (260, 480) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (260, 480) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (260, 480) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (260, 480) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (260, 480) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (260, 480) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (260, 480) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (260, 480) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (260, 480) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (260, 480) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (260, 480) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (260, 480) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (260, 480) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (260, 480) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (260, 480) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (260, 480) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (260, 480) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (260, 480) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (260, 480) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (260, 480) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (260, 480) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (260, 480) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (260, 480) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (260, 480) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (260, 480) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (260, 480) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (260, 480) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (260, 480) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (260, 480) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (260, 480) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (260, 480) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (260, 480) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (260, 480) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (260, 480) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (260, 480) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (260, 480) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (260, 480) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (260, 480) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (260, 480) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (260, 480) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (260, 480) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (260, 480) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (260, 480) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (260, 480) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (260, 480) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (260, 480) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (260, 480) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (260, 480) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (260, 480) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (260, 480) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (260, 480) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (260, 480) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (260, 480) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (260, 480) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (260, 480) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (260, 480) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (260, 480) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (260, 480) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (260, 480) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (260, 480) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (260, 480) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (260, 480) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (260, 480) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (260, 480) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (260, 480) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (260, 480) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (260, 480) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (260, 480) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (260, 480) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (260, 480) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (260, 480) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (260, 480) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (260, 480) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (260, 480) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (260, 480) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (260, 480) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (260, 480) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (260, 480) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (260, 480) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (260, 480) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (260, 480) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (260, 480) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (260, 480) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (260, 480) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (260, 480) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (260, 480) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd260;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 76
		if (frame_counter == 7'd76 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (240, 480) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (240, 480) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (240, 480) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (240, 480) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (240, 480) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (240, 480) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (240, 480) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (240, 480) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (240, 480) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (240, 480) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (240, 480) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (240, 480) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (240, 480) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (240, 480) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (240, 480) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (240, 480) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (240, 480) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (240, 480) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (240, 480) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (240, 480) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (240, 480) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (240, 480) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (240, 480) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (240, 480) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (240, 480) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (240, 480) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (240, 480) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (240, 480) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (240, 480) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (240, 480) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (240, 480) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (240, 480) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (240, 480) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (240, 480) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (240, 480) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (240, 480) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (240, 480) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (240, 480) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (240, 480) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (240, 480) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (240, 480) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (240, 480) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (240, 480) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (240, 480) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (240, 480) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (240, 480) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (240, 480) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (240, 480) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (240, 480) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (240, 480) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (240, 480) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (240, 480) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (240, 480) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (240, 480) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (240, 480) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (240, 480) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (240, 480) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (240, 480) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (240, 480) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (240, 480) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (240, 480) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (240, 480) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (240, 480) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (240, 480) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (240, 480) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (240, 480) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (240, 480) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (240, 480) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (240, 480) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (240, 480) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (240, 480) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (240, 480) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (240, 480) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (240, 480) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (240, 480) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (240, 480) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (240, 480) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (240, 480) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (240, 480) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (240, 480) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (240, 480) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (240, 480) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (240, 480) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (240, 480) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (240, 480) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (240, 480) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (240, 480) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (240, 480) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (240, 480) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (240, 480) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (240, 480) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (240, 480) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (240, 480) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (240, 480) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (240, 480) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (240, 480) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (240, 480) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (240, 480) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (240, 480) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (240, 480) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (240, 480) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (240, 480) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (240, 480) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (240, 480) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (240, 480) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (240, 480) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (240, 480) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (240, 480) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (240, 480) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (240, 480) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (240, 480) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (240, 480) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd240;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 77
		if (frame_counter == 7'd77 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (220, 480) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (220, 480) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (220, 480) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (220, 480) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (220, 480) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (220, 480) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (220, 480) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (220, 480) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (220, 480) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (220, 480) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (220, 480) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (220, 480) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (220, 480) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (220, 480) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (220, 480) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (220, 480) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (220, 480) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (220, 480) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (220, 480) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (220, 480) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (220, 480) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (220, 480) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (220, 480) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (220, 480) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (220, 480) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (220, 480) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (220, 480) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (220, 480) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (220, 480) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (220, 480) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (220, 480) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (220, 480) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (220, 480) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (220, 480) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (220, 480) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (220, 480) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (220, 480) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (220, 480) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (220, 480) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (220, 480) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (220, 480) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (220, 480) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (220, 480) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (220, 480) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (220, 480) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (220, 480) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (220, 480) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (220, 480) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (220, 480) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (220, 480) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (220, 480) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (220, 480) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (220, 480) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (220, 480) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (220, 480) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (220, 480) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (220, 480) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (220, 480) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (220, 480) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (220, 480) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (220, 480) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (220, 480) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (220, 480) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (220, 480) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (220, 480) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (220, 480) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (220, 480) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (220, 480) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (220, 480) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (220, 480) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (220, 480) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (220, 480) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (220, 480) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (220, 480) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (220, 480) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (220, 480) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (220, 480) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (220, 480) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (220, 480) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (220, 480) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (220, 480) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (220, 480) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (220, 480) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (220, 480) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (220, 480) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (220, 480) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (220, 480) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (220, 480) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (220, 480) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (220, 480) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (220, 480) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (220, 480) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (220, 480) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (220, 480) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (220, 480) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (220, 480) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (220, 480) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (220, 480) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (220, 480) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (220, 480) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (220, 480) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (220, 480) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (220, 480) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (220, 480) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (220, 480) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (220, 480) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (220, 480) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (220, 480) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (220, 480) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (220, 480) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (220, 480) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (220, 480) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd220;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 78
		if (frame_counter == 7'd78 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (200, 480) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (200, 480) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (200, 480) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (200, 480) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (200, 480) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (200, 480) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (200, 480) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (200, 480) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (200, 480) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (200, 480) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (200, 480) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (200, 480) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (200, 480) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (200, 480) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (200, 480) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (200, 480) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (200, 480) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (200, 480) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (200, 480) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (200, 480) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (200, 480) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (200, 480) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (200, 480) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (200, 480) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (200, 480) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (200, 480) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (200, 480) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (200, 480) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (200, 480) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (200, 480) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (200, 480) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (200, 480) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (200, 480) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (200, 480) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (200, 480) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (200, 480) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (200, 480) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (200, 480) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (200, 480) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (200, 480) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (200, 480) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (200, 480) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (200, 480) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (200, 480) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (200, 480) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (200, 480) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (200, 480) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (200, 480) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (200, 480) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (200, 480) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (200, 480) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (200, 480) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (200, 480) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (200, 480) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (200, 480) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (200, 480) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (200, 480) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (200, 480) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (200, 480) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (200, 480) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (200, 480) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (200, 480) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (200, 480) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (200, 480) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (200, 480) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (200, 480) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (200, 480) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (200, 480) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (200, 480) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (200, 480) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (200, 480) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (200, 480) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (200, 480) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (200, 480) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (200, 480) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (200, 480) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (200, 480) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (200, 480) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (200, 480) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (200, 480) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (200, 480) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (200, 480) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (200, 480) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (200, 480) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (200, 480) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (200, 480) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (200, 480) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (200, 480) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (200, 480) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (200, 480) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (200, 480) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (200, 480) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (200, 480) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (200, 480) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (200, 480) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (200, 480) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (200, 480) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (200, 480) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (200, 480) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (200, 480) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (200, 480) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (200, 480) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (200, 480) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (200, 480) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (200, 480) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (200, 480) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (200, 480) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (200, 480) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (200, 480) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (200, 480) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (200, 480) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (200, 480) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd200;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 79
		if (frame_counter == 7'd79 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (180, 480) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (180, 480) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (180, 480) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (180, 480) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (180, 480) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (180, 480) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (180, 480) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (180, 480) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (180, 480) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (180, 480) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (180, 480) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (180, 480) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (180, 480) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (180, 480) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (180, 480) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (180, 480) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (180, 480) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (180, 480) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (180, 480) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (180, 480) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (180, 480) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (180, 480) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (180, 480) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (180, 480) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (180, 480) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (180, 480) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (180, 480) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (180, 480) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (180, 480) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (180, 480) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (180, 480) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (180, 480) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (180, 480) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (180, 480) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (180, 480) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (180, 480) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (180, 480) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (180, 480) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (180, 480) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (180, 480) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (180, 480) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (180, 480) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (180, 480) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (180, 480) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (180, 480) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (180, 480) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (180, 480) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (180, 480) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (180, 480) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (180, 480) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (180, 480) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (180, 480) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (180, 480) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (180, 480) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (180, 480) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (180, 480) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (180, 480) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (180, 480) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (180, 480) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (180, 480) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (180, 480) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (180, 480) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (180, 480) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (180, 480) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (180, 480) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (180, 480) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (180, 480) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (180, 480) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (180, 480) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (180, 480) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (180, 480) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (180, 480) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (180, 480) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (180, 480) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (180, 480) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (180, 480) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (180, 480) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (180, 480) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (180, 480) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (180, 480) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (180, 480) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (180, 480) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (180, 480) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (180, 480) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (180, 480) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (180, 480) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (180, 480) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (180, 480) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (180, 480) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (180, 480) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (180, 480) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (180, 480) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (180, 480) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (180, 480) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (180, 480) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (180, 480) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (180, 480) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (180, 480) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (180, 480) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (180, 480) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (180, 480) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (180, 480) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (180, 480) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (180, 480) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (180, 480) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (180, 480) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (180, 480) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (180, 480) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (180, 480) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (180, 480) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (180, 480) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (180, 480) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd180;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 80
		if (frame_counter == 7'd80 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (160, 480) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (160, 480) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (160, 480) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (160, 480) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (160, 480) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (160, 480) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (160, 480) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (160, 480) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (160, 480) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (160, 480) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (160, 480) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (160, 480) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (160, 480) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (160, 480) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (160, 480) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (160, 480) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (160, 480) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (160, 480) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (160, 480) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (160, 480) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (160, 480) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (160, 480) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (160, 480) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (160, 480) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (160, 480) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (160, 480) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (160, 480) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (160, 480) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (160, 480) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (160, 480) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (160, 480) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (160, 480) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (160, 480) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (160, 480) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (160, 480) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (160, 480) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (160, 480) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (160, 480) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (160, 480) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (160, 480) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (160, 480) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (160, 480) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (160, 480) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (160, 480) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (160, 480) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (160, 480) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (160, 480) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (160, 480) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (160, 480) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (160, 480) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (160, 480) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (160, 480) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (160, 480) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (160, 480) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (160, 480) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (160, 480) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (160, 480) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (160, 480) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (160, 480) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (160, 480) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (160, 480) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (160, 480) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (160, 480) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (160, 480) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (160, 480) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (160, 480) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (160, 480) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (160, 480) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (160, 480) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (160, 480) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (160, 480) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (160, 480) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (160, 480) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (160, 480) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (160, 480) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (160, 480) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (160, 480) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (160, 480) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (160, 480) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (160, 480) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (160, 480) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (160, 480) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (160, 480) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (160, 480) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (160, 480) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (160, 480) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (160, 480) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (160, 480) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (160, 480) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (160, 480) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (160, 480) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (160, 480) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (160, 480) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (160, 480) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (160, 480) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (160, 480) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (160, 480) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (160, 480) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (160, 480) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (160, 480) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (160, 480) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (160, 480) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (160, 480) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (160, 480) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (160, 480) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (160, 480) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (160, 480) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (160, 480) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (160, 480) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (160, 480) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (160, 480) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (160, 480) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd160;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 81
		if (frame_counter == 7'd81 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (140, 480) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (140, 480) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (140, 480) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (140, 480) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (140, 480) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (140, 480) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (140, 480) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (140, 480) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (140, 480) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (140, 480) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (140, 480) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (140, 480) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (140, 480) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (140, 480) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (140, 480) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (140, 480) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (140, 480) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (140, 480) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (140, 480) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (140, 480) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (140, 480) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (140, 480) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (140, 480) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (140, 480) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (140, 480) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (140, 480) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (140, 480) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (140, 480) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (140, 480) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (140, 480) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (140, 480) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (140, 480) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (140, 480) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (140, 480) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (140, 480) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (140, 480) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (140, 480) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (140, 480) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (140, 480) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (140, 480) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (140, 480) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (140, 480) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (140, 480) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (140, 480) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (140, 480) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (140, 480) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (140, 480) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (140, 480) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (140, 480) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (140, 480) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (140, 480) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (140, 480) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (140, 480) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (140, 480) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (140, 480) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (140, 480) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (140, 480) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (140, 480) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (140, 480) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (140, 480) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (140, 480) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (140, 480) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (140, 480) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (140, 480) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (140, 480) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (140, 480) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (140, 480) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (140, 480) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (140, 480) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (140, 480) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (140, 480) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (140, 480) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (140, 480) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (140, 480) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (140, 480) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (140, 480) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (140, 480) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (140, 480) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (140, 480) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (140, 480) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (140, 480) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (140, 480) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (140, 480) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (140, 480) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (140, 480) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (140, 480) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (140, 480) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (140, 480) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (140, 480) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (140, 480) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (140, 480) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (140, 480) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (140, 480) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (140, 480) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (140, 480) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (140, 480) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (140, 480) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (140, 480) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (140, 480) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (140, 480) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (140, 480) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (140, 480) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (140, 480) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (140, 480) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (140, 480) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (140, 480) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (140, 480) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (140, 480) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (140, 480) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (140, 480) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (140, 480) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (140, 480) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd140;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 82
		if (frame_counter == 7'd82 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (120, 480) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (120, 480) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (120, 480) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (120, 480) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (120, 480) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (120, 480) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (120, 480) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (120, 480) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (120, 480) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (120, 480) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (120, 480) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (120, 480) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (120, 480) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (120, 480) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (120, 480) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (120, 480) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (120, 480) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (120, 480) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (120, 480) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (120, 480) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (120, 480) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (120, 480) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (120, 480) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (120, 480) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (120, 480) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (120, 480) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (120, 480) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (120, 480) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (120, 480) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (120, 480) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (120, 480) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (120, 480) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (120, 480) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (120, 480) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (120, 480) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (120, 480) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (120, 480) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (120, 480) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (120, 480) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (120, 480) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (120, 480) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (120, 480) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (120, 480) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (120, 480) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (120, 480) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (120, 480) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (120, 480) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (120, 480) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (120, 480) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (120, 480) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (120, 480) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (120, 480) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (120, 480) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (120, 480) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (120, 480) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (120, 480) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (120, 480) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (120, 480) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (120, 480) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (120, 480) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (120, 480) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (120, 480) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (120, 480) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (120, 480) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (120, 480) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (120, 480) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (120, 480) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (120, 480) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (120, 480) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (120, 480) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (120, 480) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (120, 480) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (120, 480) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (120, 480) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (120, 480) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (120, 480) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (120, 480) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (120, 480) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (120, 480) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (120, 480) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (120, 480) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (120, 480) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (120, 480) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (120, 480) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (120, 480) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (120, 480) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (120, 480) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (120, 480) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (120, 480) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (120, 480) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (120, 480) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (120, 480) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (120, 480) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (120, 480) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (120, 480) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (120, 480) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (120, 480) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (120, 480) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (120, 480) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (120, 480) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (120, 480) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (120, 480) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (120, 480) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (120, 480) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (120, 480) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (120, 480) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (120, 480) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (120, 480) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (120, 480) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (120, 480) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (120, 480) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (120, 480) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd120;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 83
		if (frame_counter == 7'd83 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (100, 480) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (100, 480) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (100, 480) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (100, 480) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (100, 480) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (100, 480) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (100, 480) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (100, 480) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (100, 480) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (100, 480) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (100, 480) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (100, 480) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (100, 480) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (100, 480) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (100, 480) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (100, 480) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (100, 480) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (100, 480) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (100, 480) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (100, 480) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (100, 480) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (100, 480) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (100, 480) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (100, 480) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (100, 480) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (100, 480) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (100, 480) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (100, 480) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (100, 480) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (100, 480) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (100, 480) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (100, 480) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (100, 480) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (100, 480) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (100, 480) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (100, 480) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (100, 480) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (100, 480) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (100, 480) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (100, 480) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (100, 480) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (100, 480) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (100, 480) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (100, 480) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (100, 480) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (100, 480) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (100, 480) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (100, 480) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (100, 480) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (100, 480) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (100, 480) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (100, 480) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (100, 480) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (100, 480) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (100, 480) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (100, 480) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (100, 480) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (100, 480) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (100, 480) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (100, 480) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (100, 480) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (100, 480) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (100, 480) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (100, 480) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (100, 480) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (100, 480) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (100, 480) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (100, 480) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (100, 480) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (100, 480) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (100, 480) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (100, 480) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (100, 480) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (100, 480) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (100, 480) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (100, 480) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (100, 480) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (100, 480) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (100, 480) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (100, 480) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (100, 480) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (100, 480) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (100, 480) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (100, 480) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (100, 480) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (100, 480) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (100, 480) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (100, 480) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (100, 480) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (100, 480) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (100, 480) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (100, 480) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (100, 480) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (100, 480) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (100, 480) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (100, 480) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (100, 480) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (100, 480) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (100, 480) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (100, 480) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (100, 480) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (100, 480) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (100, 480) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (100, 480) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (100, 480) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (100, 480) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (100, 480) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (100, 480) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (100, 480) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (100, 480) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (100, 480) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (100, 480) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd100;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 84
		if (frame_counter == 7'd84 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (80, 480) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (80, 480) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (80, 480) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (80, 480) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (80, 480) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (80, 480) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (80, 480) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (80, 480) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (80, 480) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (80, 480) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (80, 480) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (80, 480) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (80, 480) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (80, 480) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (80, 480) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (80, 480) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (80, 480) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (80, 480) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (80, 480) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (80, 480) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (80, 480) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (80, 480) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (80, 480) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (80, 480) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (80, 480) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (80, 480) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (80, 480) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (80, 480) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (80, 480) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (80, 480) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (80, 480) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (80, 480) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (80, 480) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (80, 480) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (80, 480) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (80, 480) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (80, 480) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (80, 480) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (80, 480) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (80, 480) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (80, 480) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (80, 480) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (80, 480) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (80, 480) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (80, 480) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (80, 480) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (80, 480) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (80, 480) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (80, 480) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (80, 480) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (80, 480) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (80, 480) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (80, 480) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (80, 480) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (80, 480) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (80, 480) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (80, 480) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (80, 480) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (80, 480) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (80, 480) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (80, 480) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (80, 480) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (80, 480) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (80, 480) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (80, 480) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (80, 480) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (80, 480) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (80, 480) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (80, 480) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (80, 480) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (80, 480) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (80, 480) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (80, 480) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (80, 480) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (80, 480) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (80, 480) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (80, 480) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (80, 480) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (80, 480) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (80, 480) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (80, 480) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (80, 480) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (80, 480) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (80, 480) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (80, 480) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (80, 480) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (80, 480) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (80, 480) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (80, 480) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (80, 480) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (80, 480) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (80, 480) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (80, 480) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (80, 480) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (80, 480) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (80, 480) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (80, 480) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (80, 480) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (80, 480) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (80, 480) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (80, 480) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (80, 480) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (80, 480) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (80, 480) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (80, 480) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (80, 480) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (80, 480) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (80, 480) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (80, 480) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (80, 480) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (80, 480) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (80, 480) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd80;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 85
		if (frame_counter == 7'd85 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (60, 480) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (60, 480) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (60, 480) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (60, 480) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (60, 480) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (60, 480) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (60, 480) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (60, 480) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (60, 480) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (60, 480) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (60, 480) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (60, 480) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (60, 480) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (60, 480) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (60, 480) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (60, 480) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (60, 480) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (60, 480) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (60, 480) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (60, 480) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (60, 480) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (60, 480) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (60, 480) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (60, 480) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (60, 480) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (60, 480) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (60, 480) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (60, 480) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (60, 480) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (60, 480) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (60, 480) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (60, 480) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (60, 480) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (60, 480) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (60, 480) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (60, 480) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (60, 480) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (60, 480) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (60, 480) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (60, 480) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (60, 480) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (60, 480) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (60, 480) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (60, 480) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (60, 480) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (60, 480) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (60, 480) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (60, 480) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (60, 480) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (60, 480) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (60, 480) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (60, 480) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (60, 480) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (60, 480) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (60, 480) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (60, 480) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (60, 480) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (60, 480) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (60, 480) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (60, 480) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (60, 480) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (60, 480) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (60, 480) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (60, 480) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (60, 480) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (60, 480) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (60, 480) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (60, 480) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (60, 480) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (60, 480) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (60, 480) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (60, 480) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (60, 480) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (60, 480) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (60, 480) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (60, 480) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (60, 480) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (60, 480) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (60, 480) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (60, 480) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (60, 480) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (60, 480) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (60, 480) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (60, 480) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (60, 480) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (60, 480) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (60, 480) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (60, 480) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (60, 480) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (60, 480) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (60, 480) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (60, 480) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (60, 480) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (60, 480) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (60, 480) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (60, 480) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (60, 480) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (60, 480) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (60, 480) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (60, 480) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (60, 480) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (60, 480) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (60, 480) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (60, 480) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (60, 480) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (60, 480) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (60, 480) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (60, 480) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (60, 480) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (60, 480) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (60, 480) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (60, 480) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd60;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 86
		if (frame_counter == 7'd86 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (40, 480) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (40, 480) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (40, 480) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (40, 480) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (40, 480) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (40, 480) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (40, 480) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (40, 480) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (40, 480) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (40, 480) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (40, 480) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (40, 480) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (40, 480) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (40, 480) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (40, 480) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (40, 480) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (40, 480) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (40, 480) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (40, 480) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (40, 480) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (40, 480) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (40, 480) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (40, 480) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (40, 480) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (40, 480) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (40, 480) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (40, 480) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (40, 480) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (40, 480) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (40, 480) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (40, 480) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (40, 480) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (40, 480) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (40, 480) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (40, 480) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (40, 480) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (40, 480) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (40, 480) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (40, 480) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (40, 480) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (40, 480) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (40, 480) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (40, 480) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (40, 480) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (40, 480) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (40, 480) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (40, 480) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (40, 480) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (40, 480) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (40, 480) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (40, 480) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (40, 480) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (40, 480) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (40, 480) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (40, 480) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (40, 480) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (40, 480) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (40, 480) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (40, 480) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (40, 480) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (40, 480) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (40, 480) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (40, 480) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (40, 480) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (40, 480) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (40, 480) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (40, 480) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (40, 480) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (40, 480) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (40, 480) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (40, 480) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (40, 480) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (40, 480) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (40, 480) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (40, 480) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (40, 480) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (40, 480) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (40, 480) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (40, 480) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (40, 480) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (40, 480) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (40, 480) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (40, 480) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (40, 480) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (40, 480) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (40, 480) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (40, 480) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (40, 480) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (40, 480) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (40, 480) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (40, 480) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (40, 480) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (40, 480) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (40, 480) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (40, 480) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (40, 480) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (40, 480) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (40, 480) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (40, 480) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (40, 480) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (40, 480) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (40, 480) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (40, 480) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (40, 480) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (40, 480) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (40, 480) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (40, 480) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (40, 480) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (40, 480) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (40, 480) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (40, 480) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (40, 480) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd40;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 87
		if (frame_counter == 7'd87 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (20, 480) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (20, 480) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (20, 480) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (20, 480) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (20, 480) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (20, 480) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (20, 480) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (20, 480) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (20, 480) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (20, 480) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (20, 480) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (20, 480) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (20, 480) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (20, 480) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (20, 480) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (20, 480) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (20, 480) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (20, 480) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (20, 480) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (20, 480) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (20, 480) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (20, 480) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (20, 480) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (20, 480) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (20, 480) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (20, 480) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (20, 480) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (20, 480) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (20, 480) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (20, 480) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (20, 480) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (20, 480) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (20, 480) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (20, 480) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (20, 480) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (20, 480) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (20, 480) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (20, 480) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (20, 480) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (20, 480) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (20, 480) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (20, 480) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (20, 480) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (20, 480) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (20, 480) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (20, 480) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (20, 480) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (20, 480) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (20, 480) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (20, 480) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (20, 480) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (20, 480) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (20, 480) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (20, 480) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (20, 480) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (20, 480) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (20, 480) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (20, 480) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (20, 480) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (20, 480) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (20, 480) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (20, 480) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (20, 480) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (20, 480) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (20, 480) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (20, 480) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (20, 480) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (20, 480) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (20, 480) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (20, 480) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (20, 480) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (20, 480) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (20, 480) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (20, 480) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (20, 480) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (20, 480) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (20, 480) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (20, 480) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (20, 480) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (20, 480) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (20, 480) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (20, 480) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (20, 480) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (20, 480) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (20, 480) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (20, 480) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (20, 480) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (20, 480) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (20, 480) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (20, 480) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (20, 480) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (20, 480) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (20, 480) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (20, 480) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (20, 480) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (20, 480) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (20, 480) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (20, 480) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (20, 480) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (20, 480) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (20, 480) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (20, 480) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (20, 480) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (20, 480) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (20, 480) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (20, 480) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (20, 480) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (20, 480) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (20, 480) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (20, 480) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (20, 480) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (20, 480) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd20;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 88
		if (frame_counter == 7'd88 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (0, 480) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (0, 480) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (0, 480) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (0, 480) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (0, 480) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (0, 480) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (0, 480) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (0, 480) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (0, 480) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (0, 480) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (0, 480) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (0, 480) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (0, 480) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (0, 480) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (0, 480) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (0, 480) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (0, 480) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (0, 480) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (0, 480) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (0, 480) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (0, 480) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (0, 480) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (0, 480) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (0, 480) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (0, 480) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (0, 480) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (0, 480) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (0, 480) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (0, 480) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (0, 480) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (0, 480) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (0, 480) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (0, 480) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (0, 480) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (0, 480) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (0, 480) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (0, 480) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (0, 480) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (0, 480) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (0, 480) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (0, 480) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (0, 480) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (0, 480) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (0, 480) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (0, 480) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (0, 480) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (0, 480) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (0, 480) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (0, 480) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (0, 480) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (0, 480) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (0, 480) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (0, 480) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (0, 480) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (0, 480) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (0, 480) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (0, 480) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (0, 480) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (0, 480) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (0, 480) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (0, 480) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (0, 480) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (0, 480) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (0, 480) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (0, 480) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (0, 480) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (0, 480) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (0, 480) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (0, 480) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (0, 480) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (0, 480) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (0, 480) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (0, 480) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (0, 480) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (0, 480) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (0, 480) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (0, 480) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (0, 480) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (0, 480) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (0, 480) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (0, 480) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (0, 480) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (0, 480) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (0, 480) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (0, 480) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (0, 480) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (0, 480) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (0, 480) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (0, 480) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (0, 480) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (0, 480) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (0, 480) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (0, 480) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (0, 480) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (0, 480) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (0, 480) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (0, 480) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (0, 480) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (0, 480) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (0, 480) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (0, 480) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (0, 480) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (0, 480) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (0, 480) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (0, 480) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (0, 480) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (0, 480) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (0, 480) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (0, 480) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (0, 480) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (0, 480) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (0, 480) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd480;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 89
		if (frame_counter == 7'd89 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (0, 460) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (0, 460) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (0, 460) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (0, 460) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (0, 460) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (0, 460) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (0, 460) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (0, 460) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (0, 460) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (0, 460) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (0, 460) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (0, 460) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (0, 460) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (0, 460) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (0, 460) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (0, 460) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (0, 460) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (0, 460) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (0, 460) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (0, 460) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (0, 460) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (0, 460) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (0, 460) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (0, 460) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (0, 460) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (0, 460) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (0, 460) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (0, 460) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (0, 460) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (0, 460) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (0, 460) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (0, 460) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (0, 460) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (0, 460) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (0, 460) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (0, 460) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (0, 460) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (0, 460) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (0, 460) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (0, 460) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (0, 460) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (0, 460) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (0, 460) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (0, 460) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (0, 460) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (0, 460) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (0, 460) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (0, 460) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (0, 460) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (0, 460) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (0, 460) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (0, 460) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (0, 460) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (0, 460) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (0, 460) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (0, 460) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (0, 460) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (0, 460) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (0, 460) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (0, 460) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (0, 460) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (0, 460) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (0, 460) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (0, 460) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (0, 460) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (0, 460) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (0, 460) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (0, 460) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (0, 460) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (0, 460) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (0, 460) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (0, 460) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (0, 460) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (0, 460) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (0, 460) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (0, 460) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (0, 460) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (0, 460) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (0, 460) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (0, 460) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (0, 460) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (0, 460) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (0, 460) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (0, 460) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (0, 460) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (0, 460) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (0, 460) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (0, 460) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (0, 460) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (0, 460) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (0, 460) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (0, 460) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (0, 460) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (0, 460) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (0, 460) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (0, 460) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (0, 460) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (0, 460) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (0, 460) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (0, 460) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (0, 460) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (0, 460) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (0, 460) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (0, 460) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (0, 460) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (0, 460) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (0, 460) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (0, 460) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (0, 460) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (0, 460) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (0, 460) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (0, 460) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd460;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 90
		if (frame_counter == 7'd90 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (0, 440) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (0, 440) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (0, 440) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (0, 440) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (0, 440) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (0, 440) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (0, 440) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (0, 440) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (0, 440) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (0, 440) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (0, 440) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (0, 440) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (0, 440) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (0, 440) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (0, 440) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (0, 440) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (0, 440) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (0, 440) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (0, 440) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (0, 440) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (0, 440) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (0, 440) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (0, 440) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (0, 440) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (0, 440) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (0, 440) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (0, 440) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (0, 440) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (0, 440) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (0, 440) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (0, 440) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (0, 440) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (0, 440) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (0, 440) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (0, 440) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (0, 440) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (0, 440) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (0, 440) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (0, 440) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (0, 440) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (0, 440) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (0, 440) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (0, 440) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (0, 440) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (0, 440) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (0, 440) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (0, 440) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (0, 440) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (0, 440) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (0, 440) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (0, 440) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (0, 440) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (0, 440) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (0, 440) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (0, 440) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (0, 440) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (0, 440) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (0, 440) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (0, 440) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (0, 440) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (0, 440) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (0, 440) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (0, 440) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (0, 440) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (0, 440) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (0, 440) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (0, 440) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (0, 440) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (0, 440) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (0, 440) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (0, 440) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (0, 440) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (0, 440) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (0, 440) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (0, 440) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (0, 440) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (0, 440) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (0, 440) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (0, 440) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (0, 440) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (0, 440) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (0, 440) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (0, 440) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (0, 440) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (0, 440) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (0, 440) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (0, 440) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (0, 440) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (0, 440) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (0, 440) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (0, 440) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (0, 440) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (0, 440) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (0, 440) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (0, 440) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (0, 440) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (0, 440) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (0, 440) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (0, 440) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (0, 440) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (0, 440) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (0, 440) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (0, 440) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (0, 440) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (0, 440) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (0, 440) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (0, 440) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (0, 440) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (0, 440) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (0, 440) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (0, 440) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (0, 440) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd440;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 91
		if (frame_counter == 7'd91 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (0, 420) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (0, 420) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (0, 420) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (0, 420) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (0, 420) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (0, 420) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (0, 420) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (0, 420) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (0, 420) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (0, 420) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (0, 420) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (0, 420) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (0, 420) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (0, 420) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (0, 420) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (0, 420) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (0, 420) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (0, 420) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (0, 420) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (0, 420) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (0, 420) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (0, 420) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (0, 420) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (0, 420) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (0, 420) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (0, 420) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (0, 420) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (0, 420) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (0, 420) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (0, 420) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (0, 420) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (0, 420) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (0, 420) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (0, 420) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (0, 420) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (0, 420) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (0, 420) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (0, 420) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (0, 420) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (0, 420) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (0, 420) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (0, 420) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (0, 420) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (0, 420) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (0, 420) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (0, 420) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (0, 420) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (0, 420) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (0, 420) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (0, 420) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (0, 420) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (0, 420) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (0, 420) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (0, 420) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (0, 420) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (0, 420) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (0, 420) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (0, 420) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (0, 420) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (0, 420) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (0, 420) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (0, 420) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (0, 420) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (0, 420) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (0, 420) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (0, 420) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (0, 420) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (0, 420) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (0, 420) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (0, 420) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (0, 420) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (0, 420) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (0, 420) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (0, 420) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (0, 420) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (0, 420) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (0, 420) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (0, 420) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (0, 420) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (0, 420) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (0, 420) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (0, 420) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (0, 420) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (0, 420) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (0, 420) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (0, 420) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (0, 420) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (0, 420) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (0, 420) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (0, 420) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (0, 420) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (0, 420) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (0, 420) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (0, 420) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (0, 420) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (0, 420) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (0, 420) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (0, 420) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (0, 420) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (0, 420) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (0, 420) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (0, 420) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (0, 420) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (0, 420) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (0, 420) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (0, 420) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (0, 420) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (0, 420) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (0, 420) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (0, 420) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (0, 420) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (0, 420) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd420;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 92
		if (frame_counter == 7'd92 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (0, 400) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (0, 400) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (0, 400) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (0, 400) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (0, 400) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (0, 400) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (0, 400) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (0, 400) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (0, 400) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (0, 400) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (0, 400) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (0, 400) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (0, 400) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (0, 400) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (0, 400) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (0, 400) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (0, 400) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (0, 400) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (0, 400) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (0, 400) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (0, 400) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (0, 400) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (0, 400) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (0, 400) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (0, 400) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (0, 400) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (0, 400) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (0, 400) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (0, 400) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (0, 400) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (0, 400) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (0, 400) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (0, 400) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (0, 400) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (0, 400) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (0, 400) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (0, 400) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (0, 400) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (0, 400) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (0, 400) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (0, 400) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (0, 400) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (0, 400) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (0, 400) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (0, 400) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (0, 400) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (0, 400) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (0, 400) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (0, 400) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (0, 400) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (0, 400) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (0, 400) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (0, 400) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (0, 400) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (0, 400) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (0, 400) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (0, 400) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (0, 400) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (0, 400) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (0, 400) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (0, 400) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (0, 400) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (0, 400) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (0, 400) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (0, 400) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (0, 400) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (0, 400) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (0, 400) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (0, 400) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (0, 400) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (0, 400) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (0, 400) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (0, 400) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (0, 400) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (0, 400) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (0, 400) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (0, 400) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (0, 400) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (0, 400) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (0, 400) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (0, 400) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (0, 400) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (0, 400) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (0, 400) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (0, 400) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (0, 400) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (0, 400) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (0, 400) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (0, 400) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (0, 400) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (0, 400) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (0, 400) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (0, 400) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (0, 400) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (0, 400) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (0, 400) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (0, 400) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (0, 400) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (0, 400) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (0, 400) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (0, 400) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (0, 400) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (0, 400) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (0, 400) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (0, 400) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (0, 400) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (0, 400) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (0, 400) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (0, 400) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (0, 400) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (0, 400) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (0, 400) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd400;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 93
		if (frame_counter == 7'd93 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (0, 380) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (0, 380) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (0, 380) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (0, 380) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (0, 380) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (0, 380) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (0, 380) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (0, 380) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (0, 380) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (0, 380) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (0, 380) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (0, 380) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (0, 380) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (0, 380) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (0, 380) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (0, 380) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (0, 380) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (0, 380) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (0, 380) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (0, 380) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (0, 380) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (0, 380) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (0, 380) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (0, 380) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (0, 380) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (0, 380) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (0, 380) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (0, 380) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (0, 380) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (0, 380) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (0, 380) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (0, 380) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (0, 380) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (0, 380) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (0, 380) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (0, 380) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (0, 380) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (0, 380) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (0, 380) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (0, 380) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (0, 380) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (0, 380) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (0, 380) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (0, 380) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (0, 380) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (0, 380) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (0, 380) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (0, 380) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (0, 380) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (0, 380) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (0, 380) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (0, 380) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (0, 380) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (0, 380) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (0, 380) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (0, 380) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (0, 380) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (0, 380) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (0, 380) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (0, 380) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (0, 380) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (0, 380) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (0, 380) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (0, 380) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (0, 380) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (0, 380) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (0, 380) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (0, 380) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (0, 380) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (0, 380) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (0, 380) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (0, 380) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (0, 380) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (0, 380) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (0, 380) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (0, 380) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (0, 380) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (0, 380) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (0, 380) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (0, 380) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (0, 380) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (0, 380) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (0, 380) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (0, 380) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (0, 380) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (0, 380) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (0, 380) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (0, 380) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (0, 380) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (0, 380) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (0, 380) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (0, 380) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (0, 380) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (0, 380) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (0, 380) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (0, 380) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (0, 380) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (0, 380) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (0, 380) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (0, 380) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (0, 380) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (0, 380) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (0, 380) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (0, 380) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (0, 380) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (0, 380) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (0, 380) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (0, 380) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (0, 380) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (0, 380) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (0, 380) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (0, 380) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd380;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 94
		if (frame_counter == 7'd94 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (0, 360) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (0, 360) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (0, 360) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (0, 360) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (0, 360) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (0, 360) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (0, 360) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (0, 360) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (0, 360) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (0, 360) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (0, 360) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (0, 360) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (0, 360) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (0, 360) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (0, 360) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (0, 360) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (0, 360) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (0, 360) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (0, 360) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (0, 360) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (0, 360) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (0, 360) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (0, 360) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (0, 360) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (0, 360) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (0, 360) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (0, 360) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (0, 360) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (0, 360) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (0, 360) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (0, 360) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (0, 360) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (0, 360) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (0, 360) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (0, 360) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (0, 360) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (0, 360) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (0, 360) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (0, 360) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (0, 360) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (0, 360) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (0, 360) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (0, 360) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (0, 360) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (0, 360) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (0, 360) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (0, 360) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (0, 360) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (0, 360) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (0, 360) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (0, 360) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (0, 360) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (0, 360) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (0, 360) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (0, 360) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (0, 360) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (0, 360) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (0, 360) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (0, 360) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (0, 360) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (0, 360) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (0, 360) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (0, 360) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (0, 360) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (0, 360) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (0, 360) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (0, 360) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (0, 360) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (0, 360) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (0, 360) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (0, 360) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (0, 360) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (0, 360) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (0, 360) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (0, 360) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (0, 360) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (0, 360) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (0, 360) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (0, 360) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (0, 360) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (0, 360) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (0, 360) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (0, 360) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (0, 360) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (0, 360) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (0, 360) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (0, 360) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (0, 360) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (0, 360) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (0, 360) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (0, 360) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (0, 360) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (0, 360) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (0, 360) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (0, 360) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (0, 360) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (0, 360) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (0, 360) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (0, 360) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (0, 360) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (0, 360) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (0, 360) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (0, 360) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (0, 360) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (0, 360) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (0, 360) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (0, 360) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (0, 360) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (0, 360) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (0, 360) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (0, 360) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (0, 360) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd360;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 95
		if (frame_counter == 7'd95 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (0, 340) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (0, 340) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (0, 340) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (0, 340) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (0, 340) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (0, 340) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (0, 340) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (0, 340) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (0, 340) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (0, 340) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (0, 340) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (0, 340) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (0, 340) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (0, 340) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (0, 340) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (0, 340) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (0, 340) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (0, 340) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (0, 340) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (0, 340) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (0, 340) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (0, 340) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (0, 340) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (0, 340) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (0, 340) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (0, 340) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (0, 340) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (0, 340) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (0, 340) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (0, 340) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (0, 340) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (0, 340) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (0, 340) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (0, 340) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (0, 340) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (0, 340) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (0, 340) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (0, 340) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (0, 340) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (0, 340) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (0, 340) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (0, 340) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (0, 340) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (0, 340) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (0, 340) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (0, 340) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (0, 340) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (0, 340) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (0, 340) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (0, 340) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (0, 340) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (0, 340) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (0, 340) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (0, 340) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (0, 340) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (0, 340) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (0, 340) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (0, 340) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (0, 340) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (0, 340) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (0, 340) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (0, 340) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (0, 340) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (0, 340) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (0, 340) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (0, 340) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (0, 340) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (0, 340) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (0, 340) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (0, 340) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (0, 340) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (0, 340) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (0, 340) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (0, 340) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (0, 340) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (0, 340) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (0, 340) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (0, 340) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (0, 340) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (0, 340) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (0, 340) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (0, 340) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (0, 340) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (0, 340) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (0, 340) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (0, 340) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (0, 340) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (0, 340) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (0, 340) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (0, 340) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (0, 340) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (0, 340) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (0, 340) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (0, 340) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (0, 340) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (0, 340) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (0, 340) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (0, 340) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (0, 340) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (0, 340) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (0, 340) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (0, 340) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (0, 340) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (0, 340) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (0, 340) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (0, 340) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (0, 340) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (0, 340) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (0, 340) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (0, 340) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (0, 340) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (0, 340) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd340;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 96
		if (frame_counter == 7'd96 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (0, 320) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (0, 320) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (0, 320) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (0, 320) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (0, 320) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (0, 320) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (0, 320) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (0, 320) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (0, 320) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (0, 320) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (0, 320) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (0, 320) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (0, 320) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (0, 320) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (0, 320) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (0, 320) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (0, 320) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (0, 320) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (0, 320) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (0, 320) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (0, 320) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (0, 320) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (0, 320) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (0, 320) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (0, 320) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (0, 320) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (0, 320) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (0, 320) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (0, 320) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (0, 320) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (0, 320) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (0, 320) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (0, 320) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (0, 320) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (0, 320) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (0, 320) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (0, 320) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (0, 320) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (0, 320) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (0, 320) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (0, 320) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (0, 320) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (0, 320) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (0, 320) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (0, 320) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (0, 320) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (0, 320) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (0, 320) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (0, 320) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (0, 320) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (0, 320) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (0, 320) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (0, 320) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (0, 320) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (0, 320) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (0, 320) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (0, 320) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (0, 320) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (0, 320) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (0, 320) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (0, 320) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (0, 320) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (0, 320) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (0, 320) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (0, 320) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (0, 320) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (0, 320) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (0, 320) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (0, 320) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (0, 320) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (0, 320) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (0, 320) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (0, 320) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (0, 320) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (0, 320) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (0, 320) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (0, 320) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (0, 320) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (0, 320) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (0, 320) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (0, 320) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (0, 320) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (0, 320) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (0, 320) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (0, 320) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (0, 320) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (0, 320) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (0, 320) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (0, 320) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (0, 320) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (0, 320) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (0, 320) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (0, 320) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (0, 320) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (0, 320) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (0, 320) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (0, 320) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (0, 320) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (0, 320) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (0, 320) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (0, 320) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (0, 320) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (0, 320) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (0, 320) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (0, 320) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (0, 320) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (0, 320) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (0, 320) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (0, 320) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (0, 320) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (0, 320) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (0, 320) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd320;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 97
		if (frame_counter == 7'd97 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (0, 300) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (0, 300) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (0, 300) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (0, 300) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (0, 300) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (0, 300) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (0, 300) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (0, 300) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (0, 300) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (0, 300) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (0, 300) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (0, 300) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (0, 300) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (0, 300) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (0, 300) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (0, 300) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (0, 300) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (0, 300) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (0, 300) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (0, 300) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (0, 300) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (0, 300) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (0, 300) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (0, 300) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (0, 300) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (0, 300) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (0, 300) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (0, 300) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (0, 300) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (0, 300) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (0, 300) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (0, 300) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (0, 300) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (0, 300) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (0, 300) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (0, 300) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (0, 300) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (0, 300) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (0, 300) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (0, 300) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (0, 300) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (0, 300) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (0, 300) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (0, 300) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (0, 300) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (0, 300) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (0, 300) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (0, 300) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (0, 300) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (0, 300) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (0, 300) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (0, 300) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (0, 300) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (0, 300) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (0, 300) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (0, 300) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (0, 300) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (0, 300) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (0, 300) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (0, 300) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (0, 300) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (0, 300) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (0, 300) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (0, 300) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (0, 300) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (0, 300) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (0, 300) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (0, 300) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (0, 300) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (0, 300) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (0, 300) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (0, 300) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (0, 300) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (0, 300) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (0, 300) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (0, 300) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (0, 300) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (0, 300) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (0, 300) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (0, 300) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (0, 300) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (0, 300) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (0, 300) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (0, 300) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (0, 300) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (0, 300) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (0, 300) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (0, 300) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (0, 300) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (0, 300) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (0, 300) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (0, 300) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (0, 300) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (0, 300) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (0, 300) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (0, 300) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (0, 300) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (0, 300) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (0, 300) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (0, 300) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (0, 300) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (0, 300) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (0, 300) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (0, 300) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (0, 300) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (0, 300) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (0, 300) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (0, 300) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (0, 300) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (0, 300) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (0, 300) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (0, 300) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd300;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 98
		if (frame_counter == 7'd98 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (0, 280) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (0, 280) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (0, 280) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (0, 280) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (0, 280) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (0, 280) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (0, 280) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (0, 280) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (0, 280) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (0, 280) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (0, 280) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (0, 280) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (0, 280) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (0, 280) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (0, 280) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (0, 280) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (0, 280) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (0, 280) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (0, 280) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (0, 280) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (0, 280) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (0, 280) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (0, 280) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (0, 280) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (0, 280) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (0, 280) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (0, 280) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (0, 280) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (0, 280) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (0, 280) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (0, 280) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (0, 280) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (0, 280) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (0, 280) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (0, 280) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (0, 280) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (0, 280) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (0, 280) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (0, 280) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (0, 280) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (0, 280) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (0, 280) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (0, 280) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (0, 280) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (0, 280) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (0, 280) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (0, 280) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (0, 280) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (0, 280) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (0, 280) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (0, 280) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (0, 280) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (0, 280) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (0, 280) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (0, 280) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (0, 280) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (0, 280) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (0, 280) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (0, 280) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (0, 280) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (0, 280) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (0, 280) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (0, 280) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (0, 280) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (0, 280) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (0, 280) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (0, 280) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (0, 280) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (0, 280) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (0, 280) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (0, 280) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (0, 280) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (0, 280) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (0, 280) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (0, 280) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (0, 280) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (0, 280) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (0, 280) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (0, 280) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (0, 280) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (0, 280) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (0, 280) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (0, 280) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (0, 280) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (0, 280) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (0, 280) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (0, 280) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (0, 280) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (0, 280) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (0, 280) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (0, 280) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (0, 280) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (0, 280) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (0, 280) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (0, 280) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (0, 280) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (0, 280) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (0, 280) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (0, 280) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (0, 280) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (0, 280) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (0, 280) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (0, 280) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (0, 280) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (0, 280) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (0, 280) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (0, 280) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (0, 280) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (0, 280) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (0, 280) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (0, 280) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (0, 280) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd280;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 99
		if (frame_counter == 7'd99 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (0, 260) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (0, 260) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (0, 260) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (0, 260) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (0, 260) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (0, 260) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (0, 260) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (0, 260) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (0, 260) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (0, 260) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (0, 260) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (0, 260) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (0, 260) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (0, 260) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (0, 260) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (0, 260) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (0, 260) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (0, 260) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (0, 260) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (0, 260) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (0, 260) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (0, 260) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (0, 260) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (0, 260) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (0, 260) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (0, 260) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (0, 260) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (0, 260) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (0, 260) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (0, 260) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (0, 260) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (0, 260) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (0, 260) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (0, 260) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (0, 260) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (0, 260) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (0, 260) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (0, 260) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (0, 260) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (0, 260) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (0, 260) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (0, 260) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (0, 260) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (0, 260) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (0, 260) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (0, 260) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (0, 260) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (0, 260) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (0, 260) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (0, 260) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (0, 260) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (0, 260) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (0, 260) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (0, 260) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (0, 260) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (0, 260) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (0, 260) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (0, 260) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (0, 260) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (0, 260) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (0, 260) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (0, 260) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (0, 260) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (0, 260) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (0, 260) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (0, 260) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (0, 260) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (0, 260) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (0, 260) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (0, 260) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (0, 260) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (0, 260) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (0, 260) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (0, 260) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (0, 260) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (0, 260) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (0, 260) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (0, 260) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (0, 260) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (0, 260) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (0, 260) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (0, 260) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (0, 260) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (0, 260) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (0, 260) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (0, 260) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (0, 260) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (0, 260) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (0, 260) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (0, 260) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (0, 260) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (0, 260) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (0, 260) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (0, 260) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (0, 260) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (0, 260) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (0, 260) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (0, 260) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (0, 260) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (0, 260) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (0, 260) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (0, 260) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (0, 260) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (0, 260) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (0, 260) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (0, 260) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (0, 260) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (0, 260) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (0, 260) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (0, 260) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (0, 260) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (0, 260) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd260;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 100
		if (frame_counter == 7'd100 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (0, 240) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (0, 240) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (0, 240) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (0, 240) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (0, 240) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (0, 240) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (0, 240) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (0, 240) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (0, 240) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (0, 240) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (0, 240) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (0, 240) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (0, 240) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (0, 240) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (0, 240) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (0, 240) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (0, 240) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (0, 240) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (0, 240) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (0, 240) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (0, 240) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (0, 240) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (0, 240) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (0, 240) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (0, 240) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (0, 240) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (0, 240) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (0, 240) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (0, 240) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (0, 240) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (0, 240) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (0, 240) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (0, 240) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (0, 240) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (0, 240) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (0, 240) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (0, 240) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (0, 240) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (0, 240) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (0, 240) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (0, 240) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (0, 240) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (0, 240) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (0, 240) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (0, 240) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (0, 240) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (0, 240) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (0, 240) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (0, 240) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (0, 240) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (0, 240) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (0, 240) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (0, 240) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (0, 240) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (0, 240) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (0, 240) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (0, 240) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (0, 240) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (0, 240) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (0, 240) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (0, 240) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (0, 240) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (0, 240) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (0, 240) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (0, 240) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (0, 240) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (0, 240) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (0, 240) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (0, 240) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (0, 240) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (0, 240) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (0, 240) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (0, 240) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (0, 240) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (0, 240) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (0, 240) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (0, 240) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (0, 240) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (0, 240) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (0, 240) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (0, 240) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (0, 240) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (0, 240) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (0, 240) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (0, 240) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (0, 240) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (0, 240) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (0, 240) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (0, 240) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (0, 240) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (0, 240) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (0, 240) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (0, 240) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (0, 240) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (0, 240) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (0, 240) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (0, 240) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (0, 240) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (0, 240) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (0, 240) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (0, 240) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (0, 240) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (0, 240) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (0, 240) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (0, 240) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (0, 240) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (0, 240) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (0, 240) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (0, 240) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (0, 240) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (0, 240) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (0, 240) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd240;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 101
		if (frame_counter == 7'd101 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (0, 220) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (0, 220) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (0, 220) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (0, 220) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (0, 220) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (0, 220) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (0, 220) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (0, 220) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (0, 220) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (0, 220) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (0, 220) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (0, 220) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (0, 220) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (0, 220) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (0, 220) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (0, 220) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (0, 220) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (0, 220) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (0, 220) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (0, 220) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (0, 220) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (0, 220) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (0, 220) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (0, 220) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (0, 220) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (0, 220) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (0, 220) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (0, 220) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (0, 220) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (0, 220) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (0, 220) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (0, 220) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (0, 220) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (0, 220) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (0, 220) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (0, 220) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (0, 220) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (0, 220) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (0, 220) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (0, 220) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (0, 220) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (0, 220) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (0, 220) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (0, 220) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (0, 220) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (0, 220) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (0, 220) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (0, 220) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (0, 220) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (0, 220) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (0, 220) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (0, 220) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (0, 220) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (0, 220) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (0, 220) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (0, 220) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (0, 220) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (0, 220) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (0, 220) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (0, 220) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (0, 220) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (0, 220) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (0, 220) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (0, 220) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (0, 220) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (0, 220) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (0, 220) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (0, 220) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (0, 220) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (0, 220) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (0, 220) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (0, 220) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (0, 220) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (0, 220) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (0, 220) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (0, 220) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (0, 220) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (0, 220) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (0, 220) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (0, 220) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (0, 220) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (0, 220) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (0, 220) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (0, 220) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (0, 220) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (0, 220) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (0, 220) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (0, 220) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (0, 220) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (0, 220) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (0, 220) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (0, 220) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (0, 220) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (0, 220) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (0, 220) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (0, 220) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (0, 220) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (0, 220) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (0, 220) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (0, 220) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (0, 220) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (0, 220) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (0, 220) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (0, 220) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (0, 220) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (0, 220) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (0, 220) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (0, 220) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (0, 220) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (0, 220) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (0, 220) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (0, 220) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd220;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 102
		if (frame_counter == 7'd102 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (0, 200) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (0, 200) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (0, 200) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (0, 200) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (0, 200) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (0, 200) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (0, 200) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (0, 200) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (0, 200) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (0, 200) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (0, 200) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (0, 200) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (0, 200) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (0, 200) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (0, 200) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (0, 200) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (0, 200) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (0, 200) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (0, 200) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (0, 200) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (0, 200) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (0, 200) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (0, 200) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (0, 200) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (0, 200) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (0, 200) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (0, 200) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (0, 200) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (0, 200) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (0, 200) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (0, 200) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (0, 200) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (0, 200) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (0, 200) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (0, 200) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (0, 200) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (0, 200) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (0, 200) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (0, 200) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (0, 200) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (0, 200) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (0, 200) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (0, 200) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (0, 200) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (0, 200) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (0, 200) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (0, 200) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (0, 200) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (0, 200) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (0, 200) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (0, 200) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (0, 200) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (0, 200) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (0, 200) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (0, 200) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (0, 200) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (0, 200) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (0, 200) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (0, 200) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (0, 200) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (0, 200) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (0, 200) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (0, 200) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (0, 200) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (0, 200) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (0, 200) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (0, 200) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (0, 200) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (0, 200) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (0, 200) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (0, 200) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (0, 200) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (0, 200) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (0, 200) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (0, 200) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (0, 200) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (0, 200) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (0, 200) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (0, 200) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (0, 200) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (0, 200) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (0, 200) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (0, 200) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (0, 200) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (0, 200) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (0, 200) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (0, 200) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (0, 200) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (0, 200) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (0, 200) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (0, 200) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (0, 200) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (0, 200) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (0, 200) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (0, 200) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (0, 200) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (0, 200) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (0, 200) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (0, 200) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (0, 200) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (0, 200) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (0, 200) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (0, 200) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (0, 200) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (0, 200) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (0, 200) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (0, 200) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (0, 200) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (0, 200) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (0, 200) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (0, 200) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (0, 200) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd200;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 103
		if (frame_counter == 7'd103 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (0, 180) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (0, 180) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (0, 180) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (0, 180) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (0, 180) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (0, 180) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (0, 180) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (0, 180) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (0, 180) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (0, 180) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (0, 180) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (0, 180) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (0, 180) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (0, 180) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (0, 180) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (0, 180) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (0, 180) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (0, 180) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (0, 180) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (0, 180) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (0, 180) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (0, 180) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (0, 180) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (0, 180) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (0, 180) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (0, 180) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (0, 180) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (0, 180) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (0, 180) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (0, 180) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (0, 180) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (0, 180) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (0, 180) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (0, 180) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (0, 180) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (0, 180) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (0, 180) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (0, 180) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (0, 180) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (0, 180) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (0, 180) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (0, 180) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (0, 180) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (0, 180) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (0, 180) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (0, 180) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (0, 180) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (0, 180) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (0, 180) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (0, 180) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (0, 180) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (0, 180) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (0, 180) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (0, 180) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (0, 180) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (0, 180) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (0, 180) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (0, 180) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (0, 180) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (0, 180) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (0, 180) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (0, 180) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (0, 180) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (0, 180) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (0, 180) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (0, 180) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (0, 180) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (0, 180) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (0, 180) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (0, 180) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (0, 180) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (0, 180) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (0, 180) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (0, 180) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (0, 180) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (0, 180) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (0, 180) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (0, 180) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (0, 180) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (0, 180) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (0, 180) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (0, 180) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (0, 180) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (0, 180) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (0, 180) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (0, 180) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (0, 180) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (0, 180) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (0, 180) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (0, 180) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (0, 180) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (0, 180) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (0, 180) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (0, 180) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (0, 180) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (0, 180) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (0, 180) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (0, 180) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (0, 180) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (0, 180) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (0, 180) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (0, 180) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (0, 180) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (0, 180) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (0, 180) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (0, 180) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (0, 180) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (0, 180) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (0, 180) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (0, 180) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (0, 180) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (0, 180) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd180;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 104
		if (frame_counter == 7'd104 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (0, 160) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (0, 160) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (0, 160) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (0, 160) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (0, 160) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (0, 160) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (0, 160) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (0, 160) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (0, 160) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (0, 160) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (0, 160) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (0, 160) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (0, 160) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (0, 160) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (0, 160) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (0, 160) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (0, 160) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (0, 160) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (0, 160) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (0, 160) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (0, 160) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (0, 160) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (0, 160) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (0, 160) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (0, 160) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (0, 160) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (0, 160) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (0, 160) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (0, 160) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (0, 160) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (0, 160) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (0, 160) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (0, 160) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (0, 160) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (0, 160) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (0, 160) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (0, 160) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (0, 160) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (0, 160) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (0, 160) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (0, 160) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (0, 160) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (0, 160) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (0, 160) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (0, 160) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (0, 160) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (0, 160) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (0, 160) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (0, 160) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (0, 160) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (0, 160) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (0, 160) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (0, 160) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (0, 160) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (0, 160) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (0, 160) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (0, 160) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (0, 160) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (0, 160) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (0, 160) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (0, 160) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (0, 160) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (0, 160) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (0, 160) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (0, 160) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (0, 160) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (0, 160) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (0, 160) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (0, 160) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (0, 160) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (0, 160) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (0, 160) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (0, 160) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (0, 160) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (0, 160) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (0, 160) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (0, 160) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (0, 160) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (0, 160) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (0, 160) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (0, 160) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (0, 160) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (0, 160) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (0, 160) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (0, 160) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (0, 160) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (0, 160) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (0, 160) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (0, 160) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (0, 160) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (0, 160) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (0, 160) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (0, 160) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (0, 160) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (0, 160) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (0, 160) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (0, 160) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (0, 160) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (0, 160) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (0, 160) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (0, 160) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (0, 160) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (0, 160) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (0, 160) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (0, 160) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (0, 160) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (0, 160) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (0, 160) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (0, 160) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (0, 160) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (0, 160) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (0, 160) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd160;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 105
		if (frame_counter == 7'd105 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (0, 140) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (0, 140) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (0, 140) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (0, 140) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (0, 140) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (0, 140) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (0, 140) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (0, 140) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (0, 140) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (0, 140) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (0, 140) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (0, 140) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (0, 140) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (0, 140) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (0, 140) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (0, 140) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (0, 140) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (0, 140) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (0, 140) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (0, 140) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (0, 140) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (0, 140) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (0, 140) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (0, 140) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (0, 140) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (0, 140) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (0, 140) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (0, 140) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (0, 140) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (0, 140) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (0, 140) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (0, 140) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (0, 140) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (0, 140) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (0, 140) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (0, 140) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (0, 140) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (0, 140) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (0, 140) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (0, 140) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (0, 140) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (0, 140) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (0, 140) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (0, 140) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (0, 140) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (0, 140) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (0, 140) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (0, 140) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (0, 140) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (0, 140) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (0, 140) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (0, 140) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (0, 140) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (0, 140) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (0, 140) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (0, 140) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (0, 140) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (0, 140) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (0, 140) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (0, 140) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (0, 140) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (0, 140) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (0, 140) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (0, 140) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (0, 140) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (0, 140) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (0, 140) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (0, 140) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (0, 140) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (0, 140) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (0, 140) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (0, 140) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (0, 140) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (0, 140) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (0, 140) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (0, 140) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (0, 140) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (0, 140) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (0, 140) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (0, 140) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (0, 140) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (0, 140) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (0, 140) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (0, 140) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (0, 140) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (0, 140) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (0, 140) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (0, 140) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (0, 140) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (0, 140) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (0, 140) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (0, 140) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (0, 140) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (0, 140) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (0, 140) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (0, 140) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (0, 140) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (0, 140) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (0, 140) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (0, 140) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (0, 140) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (0, 140) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (0, 140) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (0, 140) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (0, 140) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (0, 140) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (0, 140) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (0, 140) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (0, 140) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (0, 140) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (0, 140) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (0, 140) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd140;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 106
		if (frame_counter == 7'd106 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (0, 120) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (0, 120) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (0, 120) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (0, 120) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (0, 120) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (0, 120) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (0, 120) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (0, 120) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (0, 120) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (0, 120) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (0, 120) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (0, 120) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (0, 120) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (0, 120) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (0, 120) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (0, 120) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (0, 120) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (0, 120) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (0, 120) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (0, 120) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (0, 120) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (0, 120) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (0, 120) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (0, 120) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (0, 120) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (0, 120) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (0, 120) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (0, 120) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (0, 120) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (0, 120) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (0, 120) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (0, 120) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (0, 120) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (0, 120) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (0, 120) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (0, 120) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (0, 120) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (0, 120) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (0, 120) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (0, 120) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (0, 120) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (0, 120) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (0, 120) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (0, 120) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (0, 120) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (0, 120) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (0, 120) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (0, 120) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (0, 120) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (0, 120) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (0, 120) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (0, 120) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (0, 120) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (0, 120) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (0, 120) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (0, 120) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (0, 120) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (0, 120) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (0, 120) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (0, 120) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (0, 120) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (0, 120) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (0, 120) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (0, 120) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (0, 120) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (0, 120) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (0, 120) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (0, 120) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (0, 120) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (0, 120) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (0, 120) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (0, 120) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (0, 120) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (0, 120) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (0, 120) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (0, 120) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (0, 120) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (0, 120) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (0, 120) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (0, 120) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (0, 120) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (0, 120) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (0, 120) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (0, 120) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (0, 120) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (0, 120) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (0, 120) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (0, 120) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (0, 120) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (0, 120) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (0, 120) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (0, 120) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (0, 120) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (0, 120) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (0, 120) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (0, 120) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (0, 120) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (0, 120) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (0, 120) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (0, 120) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (0, 120) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (0, 120) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (0, 120) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (0, 120) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (0, 120) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (0, 120) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (0, 120) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (0, 120) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (0, 120) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (0, 120) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (0, 120) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (0, 120) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd120;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 107
		if (frame_counter == 7'd107 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (0, 100) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (0, 100) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (0, 100) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (0, 100) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (0, 100) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (0, 100) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (0, 100) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (0, 100) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (0, 100) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (0, 100) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (0, 100) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (0, 100) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (0, 100) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (0, 100) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (0, 100) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (0, 100) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (0, 100) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (0, 100) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (0, 100) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (0, 100) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (0, 100) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (0, 100) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (0, 100) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (0, 100) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (0, 100) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (0, 100) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (0, 100) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (0, 100) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (0, 100) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (0, 100) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (0, 100) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (0, 100) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (0, 100) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (0, 100) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (0, 100) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (0, 100) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (0, 100) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (0, 100) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (0, 100) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (0, 100) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (0, 100) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (0, 100) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (0, 100) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (0, 100) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (0, 100) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (0, 100) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (0, 100) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (0, 100) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (0, 100) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (0, 100) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (0, 100) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (0, 100) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (0, 100) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (0, 100) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (0, 100) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (0, 100) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (0, 100) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (0, 100) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (0, 100) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (0, 100) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (0, 100) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (0, 100) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (0, 100) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (0, 100) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (0, 100) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (0, 100) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (0, 100) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (0, 100) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (0, 100) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (0, 100) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (0, 100) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (0, 100) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (0, 100) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (0, 100) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (0, 100) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (0, 100) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (0, 100) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (0, 100) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (0, 100) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (0, 100) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (0, 100) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (0, 100) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (0, 100) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (0, 100) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (0, 100) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (0, 100) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (0, 100) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (0, 100) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (0, 100) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (0, 100) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (0, 100) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (0, 100) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (0, 100) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (0, 100) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (0, 100) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (0, 100) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (0, 100) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (0, 100) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (0, 100) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (0, 100) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (0, 100) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (0, 100) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (0, 100) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (0, 100) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (0, 100) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (0, 100) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (0, 100) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (0, 100) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (0, 100) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (0, 100) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (0, 100) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (0, 100) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd100;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 108
		if (frame_counter == 7'd108 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (0, 80) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (0, 80) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (0, 80) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (0, 80) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (0, 80) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (0, 80) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (0, 80) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (0, 80) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (0, 80) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (0, 80) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (0, 80) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (0, 80) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (0, 80) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (0, 80) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (0, 80) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (0, 80) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (0, 80) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (0, 80) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (0, 80) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (0, 80) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (0, 80) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (0, 80) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (0, 80) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (0, 80) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (0, 80) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (0, 80) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (0, 80) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (0, 80) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (0, 80) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (0, 80) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (0, 80) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (0, 80) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (0, 80) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (0, 80) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (0, 80) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (0, 80) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (0, 80) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (0, 80) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (0, 80) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (0, 80) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (0, 80) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (0, 80) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (0, 80) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (0, 80) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (0, 80) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (0, 80) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (0, 80) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (0, 80) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (0, 80) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (0, 80) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (0, 80) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (0, 80) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (0, 80) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (0, 80) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (0, 80) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (0, 80) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (0, 80) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (0, 80) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (0, 80) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (0, 80) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (0, 80) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (0, 80) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (0, 80) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (0, 80) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (0, 80) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (0, 80) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (0, 80) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (0, 80) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (0, 80) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (0, 80) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (0, 80) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (0, 80) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (0, 80) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (0, 80) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (0, 80) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (0, 80) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (0, 80) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (0, 80) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (0, 80) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (0, 80) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (0, 80) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (0, 80) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (0, 80) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (0, 80) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (0, 80) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (0, 80) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (0, 80) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (0, 80) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (0, 80) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (0, 80) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (0, 80) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (0, 80) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (0, 80) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (0, 80) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (0, 80) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (0, 80) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (0, 80) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (0, 80) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (0, 80) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (0, 80) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (0, 80) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (0, 80) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (0, 80) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (0, 80) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (0, 80) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (0, 80) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (0, 80) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (0, 80) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (0, 80) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (0, 80) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (0, 80) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (0, 80) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd80;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 109
		if (frame_counter == 7'd109 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (0, 60) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (0, 60) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (0, 60) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (0, 60) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (0, 60) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (0, 60) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (0, 60) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (0, 60) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (0, 60) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (0, 60) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (0, 60) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (0, 60) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (0, 60) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (0, 60) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (0, 60) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (0, 60) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (0, 60) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (0, 60) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (0, 60) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (0, 60) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (0, 60) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (0, 60) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (0, 60) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (0, 60) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (0, 60) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (0, 60) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (0, 60) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (0, 60) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (0, 60) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (0, 60) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (0, 60) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (0, 60) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (0, 60) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (0, 60) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (0, 60) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (0, 60) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (0, 60) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (0, 60) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (0, 60) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (0, 60) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (0, 60) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (0, 60) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (0, 60) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (0, 60) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (0, 60) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (0, 60) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (0, 60) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (0, 60) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (0, 60) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (0, 60) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (0, 60) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (0, 60) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (0, 60) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (0, 60) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (0, 60) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (0, 60) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (0, 60) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (0, 60) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (0, 60) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (0, 60) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (0, 60) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (0, 60) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (0, 60) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (0, 60) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (0, 60) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (0, 60) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (0, 60) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (0, 60) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (0, 60) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (0, 60) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (0, 60) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (0, 60) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (0, 60) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (0, 60) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (0, 60) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (0, 60) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (0, 60) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (0, 60) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (0, 60) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (0, 60) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (0, 60) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (0, 60) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (0, 60) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (0, 60) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (0, 60) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (0, 60) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (0, 60) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (0, 60) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (0, 60) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (0, 60) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (0, 60) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (0, 60) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (0, 60) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (0, 60) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (0, 60) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (0, 60) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (0, 60) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (0, 60) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (0, 60) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (0, 60) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (0, 60) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (0, 60) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (0, 60) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (0, 60) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (0, 60) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (0, 60) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (0, 60) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (0, 60) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (0, 60) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (0, 60) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (0, 60) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (0, 60) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd60;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 110
		if (frame_counter == 7'd110 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (0, 40) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (0, 40) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (0, 40) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (0, 40) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (0, 40) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (0, 40) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (0, 40) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (0, 40) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (0, 40) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (0, 40) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (0, 40) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (0, 40) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (0, 40) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (0, 40) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (0, 40) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (0, 40) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (0, 40) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (0, 40) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (0, 40) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (0, 40) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (0, 40) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (0, 40) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (0, 40) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (0, 40) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (0, 40) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (0, 40) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (0, 40) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (0, 40) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (0, 40) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (0, 40) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (0, 40) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (0, 40) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (0, 40) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (0, 40) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (0, 40) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (0, 40) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (0, 40) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (0, 40) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (0, 40) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (0, 40) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (0, 40) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (0, 40) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (0, 40) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (0, 40) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (0, 40) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (0, 40) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (0, 40) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (0, 40) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (0, 40) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (0, 40) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (0, 40) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (0, 40) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (0, 40) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (0, 40) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (0, 40) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (0, 40) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (0, 40) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (0, 40) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (0, 40) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (0, 40) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (0, 40) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (0, 40) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (0, 40) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (0, 40) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (0, 40) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (0, 40) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (0, 40) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (0, 40) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (0, 40) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (0, 40) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (0, 40) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (0, 40) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (0, 40) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (0, 40) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (0, 40) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (0, 40) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (0, 40) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (0, 40) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (0, 40) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (0, 40) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (0, 40) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (0, 40) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (0, 40) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (0, 40) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (0, 40) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (0, 40) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (0, 40) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (0, 40) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (0, 40) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (0, 40) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (0, 40) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (0, 40) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (0, 40) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (0, 40) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (0, 40) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (0, 40) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (0, 40) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (0, 40) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (0, 40) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (0, 40) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (0, 40) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (0, 40) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (0, 40) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (0, 40) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (0, 40) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (0, 40) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (0, 40) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (0, 40) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (0, 40) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (0, 40) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (0, 40) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (0, 40) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd40;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
		// frame 111
		if (frame_counter == 7'd111 && ~frame_complete && clear_done && ~reset && ~clear_start) begin
			color <= 1'd1;
			// line 0: (0, 20) -> (0, 0)
			if (~lines_start && lines_counter == 7'd0 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd0;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 1: (0, 20) -> (20, 0)
			if (~lines_start && lines_counter == 7'd1 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd20;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 2: (0, 20) -> (40, 0)
			if (~lines_start && lines_counter == 7'd2 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd40;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 3: (0, 20) -> (60, 0)
			if (~lines_start && lines_counter == 7'd3 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd60;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 4: (0, 20) -> (80, 0)
			if (~lines_start && lines_counter == 7'd4 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd80;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 5: (0, 20) -> (100, 0)
			if (~lines_start && lines_counter == 7'd5 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd100;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 6: (0, 20) -> (120, 0)
			if (~lines_start && lines_counter == 7'd6 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd120;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 7: (0, 20) -> (140, 0)
			if (~lines_start && lines_counter == 7'd7 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd140;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 8: (0, 20) -> (160, 0)
			if (~lines_start && lines_counter == 7'd8 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd160;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 9: (0, 20) -> (180, 0)
			if (~lines_start && lines_counter == 7'd9 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd180;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 10: (0, 20) -> (200, 0)
			if (~lines_start && lines_counter == 7'd10 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd200;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 11: (0, 20) -> (220, 0)
			if (~lines_start && lines_counter == 7'd11 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd220;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 12: (0, 20) -> (240, 0)
			if (~lines_start && lines_counter == 7'd12 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd240;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 13: (0, 20) -> (260, 0)
			if (~lines_start && lines_counter == 7'd13 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd260;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 14: (0, 20) -> (280, 0)
			if (~lines_start && lines_counter == 7'd14 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd280;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 15: (0, 20) -> (300, 0)
			if (~lines_start && lines_counter == 7'd15 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd300;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 16: (0, 20) -> (320, 0)
			if (~lines_start && lines_counter == 7'd16 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd320;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 17: (0, 20) -> (340, 0)
			if (~lines_start && lines_counter == 7'd17 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd340;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 18: (0, 20) -> (360, 0)
			if (~lines_start && lines_counter == 7'd18 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd360;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 19: (0, 20) -> (380, 0)
			if (~lines_start && lines_counter == 7'd19 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd380;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 20: (0, 20) -> (400, 0)
			if (~lines_start && lines_counter == 7'd20 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd400;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 21: (0, 20) -> (420, 0)
			if (~lines_start && lines_counter == 7'd21 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd420;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 22: (0, 20) -> (440, 0)
			if (~lines_start && lines_counter == 7'd22 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd440;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 23: (0, 20) -> (460, 0)
			if (~lines_start && lines_counter == 7'd23 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd460;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 24: (0, 20) -> (480, 0)
			if (~lines_start && lines_counter == 7'd24 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd480;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 25: (0, 20) -> (500, 0)
			if (~lines_start && lines_counter == 7'd25 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd500;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 26: (0, 20) -> (520, 0)
			if (~lines_start && lines_counter == 7'd26 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd520;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 27: (0, 20) -> (540, 0)
			if (~lines_start && lines_counter == 7'd27 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd540;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 28: (0, 20) -> (560, 0)
			if (~lines_start && lines_counter == 7'd28 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd560;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 29: (0, 20) -> (580, 0)
			if (~lines_start && lines_counter == 7'd29 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd580;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 30: (0, 20) -> (600, 0)
			if (~lines_start && lines_counter == 7'd30 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd600;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 31: (0, 20) -> (620, 0)
			if (~lines_start && lines_counter == 7'd31 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd620;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 32: (0, 20) -> (639, 0)
			if (~lines_start && lines_counter == 7'd32 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd639;
				y1 <= 11'd0;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 33: (0, 20) -> (639, 20)
			if (~lines_start && lines_counter == 7'd33 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd639;
				y1 <= 11'd20;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 34: (0, 20) -> (639, 40)
			if (~lines_start && lines_counter == 7'd34 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd639;
				y1 <= 11'd40;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 35: (0, 20) -> (639, 60)
			if (~lines_start && lines_counter == 7'd35 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd639;
				y1 <= 11'd60;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 36: (0, 20) -> (639, 80)
			if (~lines_start && lines_counter == 7'd36 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd639;
				y1 <= 11'd80;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 37: (0, 20) -> (639, 100)
			if (~lines_start && lines_counter == 7'd37 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd639;
				y1 <= 11'd100;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 38: (0, 20) -> (639, 120)
			if (~lines_start && lines_counter == 7'd38 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd639;
				y1 <= 11'd120;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 39: (0, 20) -> (639, 140)
			if (~lines_start && lines_counter == 7'd39 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd639;
				y1 <= 11'd140;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 40: (0, 20) -> (639, 160)
			if (~lines_start && lines_counter == 7'd40 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd639;
				y1 <= 11'd160;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 41: (0, 20) -> (639, 180)
			if (~lines_start && lines_counter == 7'd41 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd639;
				y1 <= 11'd180;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 42: (0, 20) -> (639, 200)
			if (~lines_start && lines_counter == 7'd42 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd639;
				y1 <= 11'd200;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 43: (0, 20) -> (639, 220)
			if (~lines_start && lines_counter == 7'd43 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd639;
				y1 <= 11'd220;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 44: (0, 20) -> (639, 240)
			if (~lines_start && lines_counter == 7'd44 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd639;
				y1 <= 11'd240;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 45: (0, 20) -> (639, 260)
			if (~lines_start && lines_counter == 7'd45 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd639;
				y1 <= 11'd260;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 46: (0, 20) -> (639, 280)
			if (~lines_start && lines_counter == 7'd46 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd639;
				y1 <= 11'd280;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 47: (0, 20) -> (639, 300)
			if (~lines_start && lines_counter == 7'd47 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd639;
				y1 <= 11'd300;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 48: (0, 20) -> (639, 320)
			if (~lines_start && lines_counter == 7'd48 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd639;
				y1 <= 11'd320;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 49: (0, 20) -> (639, 340)
			if (~lines_start && lines_counter == 7'd49 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd639;
				y1 <= 11'd340;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 50: (0, 20) -> (639, 360)
			if (~lines_start && lines_counter == 7'd50 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd639;
				y1 <= 11'd360;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 51: (0, 20) -> (639, 380)
			if (~lines_start && lines_counter == 7'd51 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd639;
				y1 <= 11'd380;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 52: (0, 20) -> (639, 400)
			if (~lines_start && lines_counter == 7'd52 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd639;
				y1 <= 11'd400;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 53: (0, 20) -> (639, 420)
			if (~lines_start && lines_counter == 7'd53 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd639;
				y1 <= 11'd420;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 54: (0, 20) -> (639, 440)
			if (~lines_start && lines_counter == 7'd54 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd639;
				y1 <= 11'd440;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 55: (0, 20) -> (639, 460)
			if (~lines_start && lines_counter == 7'd55 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd639;
				y1 <= 11'd460;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 56: (0, 20) -> (639, 479)
			if (~lines_start && lines_counter == 7'd56 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd639;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 57: (0, 20) -> (619, 479)
			if (~lines_start && lines_counter == 7'd57 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd619;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 58: (0, 20) -> (599, 479)
			if (~lines_start && lines_counter == 7'd58 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd599;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 59: (0, 20) -> (579, 479)
			if (~lines_start && lines_counter == 7'd59 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd579;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 60: (0, 20) -> (559, 479)
			if (~lines_start && lines_counter == 7'd60 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd559;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 61: (0, 20) -> (539, 479)
			if (~lines_start && lines_counter == 7'd61 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd539;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 62: (0, 20) -> (519, 479)
			if (~lines_start && lines_counter == 7'd62 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd519;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 63: (0, 20) -> (499, 479)
			if (~lines_start && lines_counter == 7'd63 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd499;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 64: (0, 20) -> (479, 479)
			if (~lines_start && lines_counter == 7'd64 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd479;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 65: (0, 20) -> (459, 479)
			if (~lines_start && lines_counter == 7'd65 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd459;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 66: (0, 20) -> (439, 479)
			if (~lines_start && lines_counter == 7'd66 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd439;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 67: (0, 20) -> (419, 479)
			if (~lines_start && lines_counter == 7'd67 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd419;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 68: (0, 20) -> (399, 479)
			if (~lines_start && lines_counter == 7'd68 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd399;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 69: (0, 20) -> (379, 479)
			if (~lines_start && lines_counter == 7'd69 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd379;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 70: (0, 20) -> (359, 479)
			if (~lines_start && lines_counter == 7'd70 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd359;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 71: (0, 20) -> (339, 479)
			if (~lines_start && lines_counter == 7'd71 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd339;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 72: (0, 20) -> (319, 479)
			if (~lines_start && lines_counter == 7'd72 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd319;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 73: (0, 20) -> (299, 479)
			if (~lines_start && lines_counter == 7'd73 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd299;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 74: (0, 20) -> (279, 479)
			if (~lines_start && lines_counter == 7'd74 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd279;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 75: (0, 20) -> (259, 479)
			if (~lines_start && lines_counter == 7'd75 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd259;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 76: (0, 20) -> (239, 479)
			if (~lines_start && lines_counter == 7'd76 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd239;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 77: (0, 20) -> (219, 479)
			if (~lines_start && lines_counter == 7'd77 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd219;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 78: (0, 20) -> (199, 479)
			if (~lines_start && lines_counter == 7'd78 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd199;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 79: (0, 20) -> (179, 479)
			if (~lines_start && lines_counter == 7'd79 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd179;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 80: (0, 20) -> (159, 479)
			if (~lines_start && lines_counter == 7'd80 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd159;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 81: (0, 20) -> (139, 479)
			if (~lines_start && lines_counter == 7'd81 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd139;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 82: (0, 20) -> (119, 479)
			if (~lines_start && lines_counter == 7'd82 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd119;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 83: (0, 20) -> (99, 479)
			if (~lines_start && lines_counter == 7'd83 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd99;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 84: (0, 20) -> (79, 479)
			if (~lines_start && lines_counter == 7'd84 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd79;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 85: (0, 20) -> (59, 479)
			if (~lines_start && lines_counter == 7'd85 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd59;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 86: (0, 20) -> (39, 479)
			if (~lines_start && lines_counter == 7'd86 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd39;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 87: (0, 20) -> (19, 479)
			if (~lines_start && lines_counter == 7'd87 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd19;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 88: (0, 20) -> (0, 479)
			if (~lines_start && lines_counter == 7'd88 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd0;
				y1 <= 11'd479;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 89: (0, 20) -> (0, 459)
			if (~lines_start && lines_counter == 7'd89 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd0;
				y1 <= 11'd459;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 90: (0, 20) -> (0, 439)
			if (~lines_start && lines_counter == 7'd90 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd0;
				y1 <= 11'd439;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 91: (0, 20) -> (0, 419)
			if (~lines_start && lines_counter == 7'd91 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd0;
				y1 <= 11'd419;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 92: (0, 20) -> (0, 399)
			if (~lines_start && lines_counter == 7'd92 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd0;
				y1 <= 11'd399;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 93: (0, 20) -> (0, 379)
			if (~lines_start && lines_counter == 7'd93 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd0;
				y1 <= 11'd379;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 94: (0, 20) -> (0, 359)
			if (~lines_start && lines_counter == 7'd94 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd0;
				y1 <= 11'd359;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 95: (0, 20) -> (0, 339)
			if (~lines_start && lines_counter == 7'd95 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd0;
				y1 <= 11'd339;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 96: (0, 20) -> (0, 319)
			if (~lines_start && lines_counter == 7'd96 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd0;
				y1 <= 11'd319;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 97: (0, 20) -> (0, 299)
			if (~lines_start && lines_counter == 7'd97 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd0;
				y1 <= 11'd299;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 98: (0, 20) -> (0, 279)
			if (~lines_start && lines_counter == 7'd98 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd0;
				y1 <= 11'd279;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 99: (0, 20) -> (0, 259)
			if (~lines_start && lines_counter == 7'd99 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd0;
				y1 <= 11'd259;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 100: (0, 20) -> (0, 239)
			if (~lines_start && lines_counter == 7'd100 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd0;
				y1 <= 11'd239;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 101: (0, 20) -> (0, 219)
			if (~lines_start && lines_counter == 7'd101 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd0;
				y1 <= 11'd219;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 102: (0, 20) -> (0, 199)
			if (~lines_start && lines_counter == 7'd102 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd0;
				y1 <= 11'd199;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 103: (0, 20) -> (0, 179)
			if (~lines_start && lines_counter == 7'd103 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd0;
				y1 <= 11'd179;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 104: (0, 20) -> (0, 159)
			if (~lines_start && lines_counter == 7'd104 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd0;
				y1 <= 11'd159;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 105: (0, 20) -> (0, 139)
			if (~lines_start && lines_counter == 7'd105 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd0;
				y1 <= 11'd139;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 106: (0, 20) -> (0, 119)
			if (~lines_start && lines_counter == 7'd106 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd0;
				y1 <= 11'd119;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 107: (0, 20) -> (0, 99)
			if (~lines_start && lines_counter == 7'd107 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd0;
				y1 <= 11'd99;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 108: (0, 20) -> (0, 79)
			if (~lines_start && lines_counter == 7'd108 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd0;
				y1 <= 11'd79;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 109: (0, 20) -> (0, 59)
			if (~lines_start && lines_counter == 7'd109 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd0;
				y1 <= 11'd59;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 110: (0, 20) -> (0, 39)
			if (~lines_start && lines_counter == 7'd110 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd0;
				y1 <= 11'd39;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
			end
			// line 111: (0, 20) -> (0, 19)
			if (~lines_start && lines_counter == 7'd111 && lines_done) begin
				x0 <= 11'd0;
				y0 <= 11'd20;
				x1 <= 11'd0;
				y1 <= 11'd19;
				lines_start <= 1'd1;
				lines_counter <= lines_counter + 1'd1;
				//frame is complete
				lines_counter <= 7'd0;
				frame_complete <= 1'd1;
			end
		end
	end
endmodule // fancy_animation


module fancy_animation_testbench();
    logic clk, reset;
    logic done, color;
    logic [10:0] x, y;

fancy_animation dut(.*);

    // simulated clock
	parameter period = 100;
    initial begin
        clk <= 0;
        forever begin
            #(period/2)
            clk <= ~clk;
        end
    end

    // begin tests
	initial begin
        // Pre-test setup
        reset <= 1; repeat(500) @(posedge clk);
        // Test 1: animation
        // Expected: x, y should iterate through all coordinates of the VGA signal,
        //           and clears itself repeatedly.
		reset <= 0; repeat(5000) @(posedge clk);        // Test 2: clear screen
        reset <= 1; repeat(500) @(posedge clk);
        $stop;
    end

endmodule // fancy_animation_testbench
